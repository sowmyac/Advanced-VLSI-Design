*
*
*
*                       LINUX           Thu Jul  3 17:34:39 2014
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - QRC - (32-bit)
*  Version        : 9.1.3-p005
*  Build Date     : Tue Aug  3 12:36:00 PDT 2010
*
*  HSPICE LIBRARY
*
*
*
*.GLOBAL vdd vss
*
.SUBCKT SRAM vdd vss wr clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 addr_en data0 data1
+ data2 data3 data4 data5 data6 data7 data8 data9
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MI0/I4060/T2	BL36	net955	I0/I4060/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4052/T2	BL36	net954	I0/I4052/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4051/T2	BL36	net953	I0/I4051/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4076/T2	BL36	net952	I0/I4076/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4057/T2	BL36	net951	I0/I4057/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4072/T2	BL36	net950	I0/I4072/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4070/T2	BL36	net949	I0/I4070/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4066/T2	BL36	net948	I0/I4066/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4058/T2	BL36	net947	I0/I4058/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4060/T5	I0/I4060/net13	I0/I4060/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4052/T5	I0/I4052/net13	I0/I4052/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4051/T5	I0/I4051/net13	I0/I4051/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4076/T5	I0/I4076/net13	I0/I4076/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4057/T5	I0/I4057/net13	I0/I4057/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4072/T5	I0/I4072/net13	I0/I4072/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4070/T5	I0/I4070/net13	I0/I4070/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4066/T5	I0/I4066/net13	I0/I4066/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4058/T5	I0/I4058/net13	I0/I4058/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4060/T4	vss	I0/I4060/net13	I0/I4060/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4052/T4	vss	I0/I4052/net13	I0/I4052/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4051/T4	vss	I0/I4051/net13	I0/I4051/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4076/T4	vss	I0/I4076/net13	I0/I4076/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4057/T4	vss	I0/I4057/net13	I0/I4057/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4072/T4	vss	I0/I4072/net13	I0/I4072/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4070/T4	vss	I0/I4070/net13	I0/I4070/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4066/T4	vss	I0/I4066/net13	I0/I4066/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4058/T4	vss	I0/I4058/net13	I0/I4058/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4060/T3	I0/I4060/net049	net955	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4052/T3	I0/I4052/net049	net954	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4051/T3	I0/I4051/net049	net953	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4076/T3	I0/I4076/net049	net952	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4057/T3	I0/I4057/net049	net951	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4072/T3	I0/I4072/net049	net950	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4070/T3	I0/I4070/net049	net949	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4066/T3	I0/I4066/net049	net948	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4058/T3	I0/I4058/net049	net947	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4156/T4	vss	I0/I4156/net13	I0/I4156/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4148/T4	vss	I0/I4148/net13	I0/I4148/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4156/T5	I0/I4156/net13	I0/I4156/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4148/T5	I0/I4148/net13	I0/I4148/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4156/T2	BL37	net955	I0/I4156/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4148/T2	BL37	net954	I0/I4148/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4147/T4	vss	I0/I4147/net13	I0/I4147/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4172/T4	vss	I0/I4172/net13	I0/I4172/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4147/T5	I0/I4147/net13	I0/I4147/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4172/T5	I0/I4172/net13	I0/I4172/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4147/T2	BL37	net953	I0/I4147/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4172/T2	BL37	net952	I0/I4172/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4153/T4	vss	I0/I4153/net13	I0/I4153/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4153/T5	I0/I4153/net13	I0/I4153/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4153/T2	BL37	net951	I0/I4153/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4168/T4	vss	I0/I4168/net13	I0/I4168/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4166/T4	vss	I0/I4166/net13	I0/I4166/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4168/T5	I0/I4168/net13	I0/I4168/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4166/T5	I0/I4166/net13	I0/I4166/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4168/T2	BL37	net950	I0/I4168/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4166/T2	BL37	net949	I0/I4166/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4162/T4	vss	I0/I4162/net13	I0/I4162/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4154/T4	vss	I0/I4154/net13	I0/I4154/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4162/T5	I0/I4162/net13	I0/I4162/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4154/T5	I0/I4154/net13	I0/I4154/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4162/T2	BL37	net948	I0/I4162/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4154/T2	BL37	net947	I0/I4154/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4156/T3	I0/I4156/net049	net955	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4148/T3	I0/I4148/net049	net954	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4147/T3	I0/I4147/net049	net953	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4172/T3	I0/I4172/net049	net952	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4153/T3	I0/I4153/net049	net951	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4168/T3	I0/I4168/net049	net950	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4166/T3	I0/I4166/net049	net949	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4162/T3	I0/I4162/net049	net948	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4154/T3	I0/I4154/net049	net947	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4220/T5	I0/I4220/net13	I0/I4220/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4220/T2	BL39	net955	I0/I4220/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4188/T3	I0/I4188/net049	net955	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4188/T4	vss	I0/I4188/net13	I0/I4188/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4188/T5	I0/I4188/net13	I0/I4188/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4188/T2	BL38	net955	I0/I4188/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4212/T5	I0/I4212/net13	I0/I4212/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4212/T2	BL39	net954	I0/I4212/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4180/T3	I0/I4180/net049	net954	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4180/T4	vss	I0/I4180/net13	I0/I4180/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4180/T5	I0/I4180/net13	I0/I4180/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4180/T2	BL38	net954	I0/I4180/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4211/T5	I0/I4211/net13	I0/I4211/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4211/T2	BL39	net953	I0/I4211/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4179/T3	I0/I4179/net049	net953	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4179/T4	vss	I0/I4179/net13	I0/I4179/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4179/T5	I0/I4179/net13	I0/I4179/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4179/T2	BL38	net953	I0/I4179/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4236/T5	I0/I4236/net13	I0/I4236/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4236/T2	BL39	net952	I0/I4236/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4204/T3	I0/I4204/net049	net952	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4204/T4	vss	I0/I4204/net13	I0/I4204/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4204/T5	I0/I4204/net13	I0/I4204/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4204/T2	BL38	net952	I0/I4204/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4217/T5	I0/I4217/net13	I0/I4217/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4217/T2	BL39	net951	I0/I4217/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4185/T3	I0/I4185/net049	net951	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4185/T4	vss	I0/I4185/net13	I0/I4185/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4185/T5	I0/I4185/net13	I0/I4185/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4185/T2	BL38	net951	I0/I4185/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4232/T5	I0/I4232/net13	I0/I4232/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4232/T2	BL39	net950	I0/I4232/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4200/T3	I0/I4200/net049	net950	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4200/T4	vss	I0/I4200/net13	I0/I4200/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4200/T5	I0/I4200/net13	I0/I4200/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4200/T2	BL38	net950	I0/I4200/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4230/T5	I0/I4230/net13	I0/I4230/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4230/T2	BL39	net949	I0/I4230/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4198/T3	I0/I4198/net049	net949	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4198/T4	vss	I0/I4198/net13	I0/I4198/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4198/T5	I0/I4198/net13	I0/I4198/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4198/T2	BL38	net949	I0/I4198/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4226/T5	I0/I4226/net13	I0/I4226/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4226/T2	BL39	net948	I0/I4226/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4194/T3	I0/I4194/net049	net948	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4194/T4	vss	I0/I4194/net13	I0/I4194/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4194/T5	I0/I4194/net13	I0/I4194/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4194/T2	BL38	net948	I0/I4194/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4218/T5	I0/I4218/net13	I0/I4218/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4218/T2	BL39	net947	I0/I4218/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4186/T3	I0/I4186/net049	net947	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4186/T4	vss	I0/I4186/net13	I0/I4186/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4186/T5	I0/I4186/net13	I0/I4186/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4186/T2	BL38	net947	I0/I4186/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4059/T2	BL36	net946	I0/I4059/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4049/T2	BL36	net945	I0/I4049/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4075/T2	BL36	net944	I0/I4075/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4069/T2	BL36	net943	I0/I4069/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4055/T2	BL36	net942	I0/I4055/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4048/T2	BL36	net941	I0/I4048/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4071/T2	BL36	net940	I0/I4071/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4068/T2	BL36	net939	I0/I4068/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4046/T2	BL36	net938	I0/I4046/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4059/T5	I0/I4059/net13	I0/I4059/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4049/T5	I0/I4049/net13	I0/I4049/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4075/T5	I0/I4075/net13	I0/I4075/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4069/T5	I0/I4069/net13	I0/I4069/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4055/T5	I0/I4055/net13	I0/I4055/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4048/T5	I0/I4048/net13	I0/I4048/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4071/T5	I0/I4071/net13	I0/I4071/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4068/T5	I0/I4068/net13	I0/I4068/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4046/T5	I0/I4046/net13	I0/I4046/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4059/T4	vss	I0/I4059/net13	I0/I4059/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4049/T4	vss	I0/I4049/net13	I0/I4049/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4075/T4	vss	I0/I4075/net13	I0/I4075/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4069/T4	vss	I0/I4069/net13	I0/I4069/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4055/T4	vss	I0/I4055/net13	I0/I4055/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4048/T4	vss	I0/I4048/net13	I0/I4048/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4071/T4	vss	I0/I4071/net13	I0/I4071/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4068/T4	vss	I0/I4068/net13	I0/I4068/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4046/T4	vss	I0/I4046/net13	I0/I4046/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4059/T3	I0/I4059/net049	net946	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4049/T3	I0/I4049/net049	net945	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4075/T3	I0/I4075/net049	net944	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4069/T3	I0/I4069/net049	net943	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4055/T3	I0/I4055/net049	net942	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4048/T3	I0/I4048/net049	net941	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4071/T3	I0/I4071/net049	net940	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4068/T3	I0/I4068/net049	net939	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4046/T3	I0/I4046/net049	net938	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4155/T4	vss	I0/I4155/net13	I0/I4155/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4145/T4	vss	I0/I4145/net13	I0/I4145/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4155/T5	I0/I4155/net13	I0/I4155/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4145/T5	I0/I4145/net13	I0/I4145/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4155/T2	BL37	net946	I0/I4155/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4145/T2	BL37	net945	I0/I4145/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4171/T4	vss	I0/I4171/net13	I0/I4171/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4165/T4	vss	I0/I4165/net13	I0/I4165/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4171/T5	I0/I4171/net13	I0/I4171/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4165/T5	I0/I4165/net13	I0/I4165/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4171/T2	BL37	net944	I0/I4171/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4165/T2	BL37	net943	I0/I4165/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4151/T4	vss	I0/I4151/net13	I0/I4151/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4151/T5	I0/I4151/net13	I0/I4151/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4151/T2	BL37	net942	I0/I4151/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4144/T4	vss	I0/I4144/net13	I0/I4144/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4167/T4	vss	I0/I4167/net13	I0/I4167/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4144/T5	I0/I4144/net13	I0/I4144/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4167/T5	I0/I4167/net13	I0/I4167/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4144/T2	BL37	net941	I0/I4144/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4167/T2	BL37	net940	I0/I4167/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4164/T4	vss	I0/I4164/net13	I0/I4164/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4142/T4	vss	I0/I4142/net13	I0/I4142/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4164/T5	I0/I4164/net13	I0/I4164/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4142/T5	I0/I4142/net13	I0/I4142/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4164/T2	BL37	net939	I0/I4164/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4142/T2	BL37	net938	I0/I4142/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4155/T3	I0/I4155/net049	net946	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4145/T3	I0/I4145/net049	net945	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4171/T3	I0/I4171/net049	net944	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4165/T3	I0/I4165/net049	net943	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4151/T3	I0/I4151/net049	net942	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4144/T3	I0/I4144/net049	net941	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4167/T3	I0/I4167/net049	net940	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4164/T3	I0/I4164/net049	net939	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4142/T3	I0/I4142/net049	net938	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4219/T5	I0/I4219/net13	I0/I4219/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4219/T2	BL39	net946	I0/I4219/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4187/T3	I0/I4187/net049	net946	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4187/T4	vss	I0/I4187/net13	I0/I4187/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4187/T5	I0/I4187/net13	I0/I4187/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4187/T2	BL38	net946	I0/I4187/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4209/T5	I0/I4209/net13	I0/I4209/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4209/T2	BL39	net945	I0/I4209/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4177/T3	I0/I4177/net049	net945	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4177/T4	vss	I0/I4177/net13	I0/I4177/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4177/T5	I0/I4177/net13	I0/I4177/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4177/T2	BL38	net945	I0/I4177/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4235/T5	I0/I4235/net13	I0/I4235/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4235/T2	BL39	net944	I0/I4235/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4203/T3	I0/I4203/net049	net944	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4203/T4	vss	I0/I4203/net13	I0/I4203/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4203/T5	I0/I4203/net13	I0/I4203/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4203/T2	BL38	net944	I0/I4203/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4229/T5	I0/I4229/net13	I0/I4229/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4229/T2	BL39	net943	I0/I4229/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4197/T3	I0/I4197/net049	net943	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4197/T4	vss	I0/I4197/net13	I0/I4197/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4197/T5	I0/I4197/net13	I0/I4197/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4197/T2	BL38	net943	I0/I4197/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4215/T5	I0/I4215/net13	I0/I4215/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4215/T2	BL39	net942	I0/I4215/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4183/T3	I0/I4183/net049	net942	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4183/T4	vss	I0/I4183/net13	I0/I4183/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4183/T5	I0/I4183/net13	I0/I4183/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4183/T2	BL38	net942	I0/I4183/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4208/T5	I0/I4208/net13	I0/I4208/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4208/T2	BL39	net941	I0/I4208/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4176/T3	I0/I4176/net049	net941	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4176/T4	vss	I0/I4176/net13	I0/I4176/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4176/T5	I0/I4176/net13	I0/I4176/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4176/T2	BL38	net941	I0/I4176/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4231/T5	I0/I4231/net13	I0/I4231/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4231/T2	BL39	net940	I0/I4231/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4199/T3	I0/I4199/net049	net940	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4199/T4	vss	I0/I4199/net13	I0/I4199/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4199/T5	I0/I4199/net13	I0/I4199/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4199/T2	BL38	net940	I0/I4199/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4228/T5	I0/I4228/net13	I0/I4228/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4228/T2	BL39	net939	I0/I4228/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4196/T3	I0/I4196/net049	net939	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4196/T4	vss	I0/I4196/net13	I0/I4196/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4196/T5	I0/I4196/net13	I0/I4196/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4196/T2	BL38	net939	I0/I4196/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4206/T5	I0/I4206/net13	I0/I4206/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4206/T2	BL39	net938	I0/I4206/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4174/T3	I0/I4174/net049	net938	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4174/T4	vss	I0/I4174/net13	I0/I4174/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4174/T5	I0/I4174/net13	I0/I4174/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4174/T2	BL38	net938	I0/I4174/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4143/T4	vss	I0/I4143/net13	I0/I4143/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4143/T5	I0/I4143/net13	I0/I4143/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4143/T2	BL37	net937	I0/I4143/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4047/T3	I0/I4047/net049	net937	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4047/T4	vss	I0/I4047/net13	I0/I4047/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4047/T5	I0/I4047/net13	I0/I4047/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4047/T2	BL36	net937	I0/I4047/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4143/T3	I0/I4143/net049	net937	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4207/T5	I0/I4207/net13	I0/I4207/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4207/T2	BL39	net937	I0/I4207/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4175/T3	I0/I4175/net049	net937	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4175/T4	vss	I0/I4175/net13	I0/I4175/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4175/T5	I0/I4175/net13	I0/I4175/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4175/T2	BL38	net937	I0/I4175/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4150/T4	vss	I0/I4150/net13	I0/I4150/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4150/T5	I0/I4150/net13	I0/I4150/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4150/T2	BL37	net936	I0/I4150/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4054/T3	I0/I4054/net049	net936	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4054/T4	vss	I0/I4054/net13	I0/I4054/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4054/T5	I0/I4054/net13	I0/I4054/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4054/T2	BL36	net936	I0/I4054/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4150/T3	I0/I4150/net049	net936	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4214/T5	I0/I4214/net13	I0/I4214/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4214/T2	BL39	net936	I0/I4214/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4182/T3	I0/I4182/net049	net936	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4182/T4	vss	I0/I4182/net13	I0/I4182/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4182/T5	I0/I4182/net13	I0/I4182/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4182/T2	BL38	net936	I0/I4182/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4152/T4	vss	I0/I4152/net13	I0/I4152/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4152/T5	I0/I4152/net13	I0/I4152/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4152/T2	BL37	net935	I0/I4152/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4056/T3	I0/I4056/net049	net935	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4056/T4	vss	I0/I4056/net13	I0/I4056/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4056/T5	I0/I4056/net13	I0/I4056/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4056/T2	BL36	net935	I0/I4056/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4152/T3	I0/I4152/net049	net935	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4216/T5	I0/I4216/net13	I0/I4216/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4216/T2	BL39	net935	I0/I4216/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4184/T3	I0/I4184/net049	net935	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4184/T4	vss	I0/I4184/net13	I0/I4184/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4184/T5	I0/I4184/net13	I0/I4184/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4184/T2	BL38	net935	I0/I4184/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4158/T4	vss	I0/I4158/net13	I0/I4158/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4158/T5	I0/I4158/net13	I0/I4158/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4158/T2	BL37	net934	I0/I4158/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4062/T3	I0/I4062/net049	net934	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4062/T4	vss	I0/I4062/net13	I0/I4062/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4062/T5	I0/I4062/net13	I0/I4062/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4062/T2	BL36	net934	I0/I4062/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4158/T3	I0/I4158/net049	net934	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4222/T5	I0/I4222/net13	I0/I4222/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4222/T2	BL39	net934	I0/I4222/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4190/T3	I0/I4190/net049	net934	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4190/T4	vss	I0/I4190/net13	I0/I4190/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4190/T5	I0/I4190/net13	I0/I4190/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4190/T2	BL38	net934	I0/I4190/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4160/T4	vss	I0/I4160/net13	I0/I4160/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4160/T5	I0/I4160/net13	I0/I4160/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4160/T2	BL37	net933	I0/I4160/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4064/T3	I0/I4064/net049	net933	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4064/T4	vss	I0/I4064/net13	I0/I4064/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4064/T5	I0/I4064/net13	I0/I4064/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4064/T2	BL36	net933	I0/I4064/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4160/T3	I0/I4160/net049	net933	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4224/T5	I0/I4224/net13	I0/I4224/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4224/T2	BL39	net933	I0/I4224/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4192/T3	I0/I4192/net049	net933	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4192/T4	vss	I0/I4192/net13	I0/I4192/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4192/T5	I0/I4192/net13	I0/I4192/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4192/T2	BL38	net933	I0/I4192/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4149/T4	vss	I0/I4149/net13	I0/I4149/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4149/T5	I0/I4149/net13	I0/I4149/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4149/T2	BL37	net932	I0/I4149/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4053/T3	I0/I4053/net049	net932	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4053/T4	vss	I0/I4053/net13	I0/I4053/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4053/T5	I0/I4053/net13	I0/I4053/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4053/T2	BL36	net932	I0/I4053/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4149/T3	I0/I4149/net049	net932	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4213/T5	I0/I4213/net13	I0/I4213/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4213/T2	BL39	net932	I0/I4213/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4181/T3	I0/I4181/net049	net932	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4181/T4	vss	I0/I4181/net13	I0/I4181/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4181/T5	I0/I4181/net13	I0/I4181/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4181/T2	BL38	net932	I0/I4181/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4163/T4	vss	I0/I4163/net13	I0/I4163/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4163/T5	I0/I4163/net13	I0/I4163/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4163/T2	BL37	net931	I0/I4163/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4067/T3	I0/I4067/net049	net931	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4067/T4	vss	I0/I4067/net13	I0/I4067/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4067/T5	I0/I4067/net13	I0/I4067/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4067/T2	BL36	net931	I0/I4067/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4163/T3	I0/I4163/net049	net931	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4227/T5	I0/I4227/net13	I0/I4227/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4227/T2	BL39	net931	I0/I4227/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4195/T3	I0/I4195/net049	net931	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4195/T4	vss	I0/I4195/net13	I0/I4195/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4195/T5	I0/I4195/net13	I0/I4195/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4195/T2	BL38	net931	I0/I4195/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4157/T4	vss	I0/I4157/net13	I0/I4157/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4157/T5	I0/I4157/net13	I0/I4157/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4157/T2	BL37	net930	I0/I4157/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4061/T3	I0/I4061/net049	net930	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4061/T4	vss	I0/I4061/net13	I0/I4061/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4061/T5	I0/I4061/net13	I0/I4061/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4061/T2	BL36	net930	I0/I4061/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4157/T3	I0/I4157/net049	net930	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4221/T5	I0/I4221/net13	I0/I4221/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4221/T2	BL39	net930	I0/I4221/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4189/T3	I0/I4189/net049	net930	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4189/T4	vss	I0/I4189/net13	I0/I4189/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4189/T5	I0/I4189/net13	I0/I4189/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4189/T2	BL38	net930	I0/I4189/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4161/T4	vss	I0/I4161/net13	I0/I4161/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4161/T5	I0/I4161/net13	I0/I4161/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4161/T2	BL37	net929	I0/I4161/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4065/T3	I0/I4065/net049	net929	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4065/T4	vss	I0/I4065/net13	I0/I4065/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4065/T5	I0/I4065/net13	I0/I4065/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4065/T2	BL36	net929	I0/I4065/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4161/T3	I0/I4161/net049	net929	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4225/T5	I0/I4225/net13	I0/I4225/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4225/T2	BL39	net929	I0/I4225/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4193/T3	I0/I4193/net049	net929	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4193/T4	vss	I0/I4193/net13	I0/I4193/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4193/T5	I0/I4193/net13	I0/I4193/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4193/T2	BL38	net929	I0/I4193/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4173/T4	vss	I0/I4173/net13	I0/I4173/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4173/T5	I0/I4173/net13	I0/I4173/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4173/T2	BL37	net928	I0/I4173/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4077/T3	I0/I4077/net049	net928	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4077/T4	vss	I0/I4077/net13	I0/I4077/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4077/T5	I0/I4077/net13	I0/I4077/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4077/T2	BL36	net928	I0/I4077/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4173/T3	I0/I4173/net049	net928	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4237/T5	I0/I4237/net13	I0/I4237/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4237/T2	BL39	net928	I0/I4237/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4205/T3	I0/I4205/net049	net928	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4205/T4	vss	I0/I4205/net13	I0/I4205/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4205/T5	I0/I4205/net13	I0/I4205/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4205/T2	BL38	net928	I0/I4205/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4159/T4	vss	I0/I4159/net13	I0/I4159/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4159/T5	I0/I4159/net13	I0/I4159/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4159/T2	BL37	net927	I0/I4159/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4063/T3	I0/I4063/net049	net927	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4063/T4	vss	I0/I4063/net13	I0/I4063/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4063/T5	I0/I4063/net13	I0/I4063/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4063/T2	BL36	net927	I0/I4063/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4159/T3	I0/I4159/net049	net927	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4223/T5	I0/I4223/net13	I0/I4223/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4223/T2	BL39	net927	I0/I4223/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4191/T3	I0/I4191/net049	net927	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4191/T4	vss	I0/I4191/net13	I0/I4191/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4191/T5	I0/I4191/net13	I0/I4191/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4191/T2	BL38	net927	I0/I4191/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4170/T4	vss	I0/I4170/net13	I0/I4170/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4170/T5	I0/I4170/net13	I0/I4170/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4170/T2	BL37	net926	I0/I4170/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4074/T3	I0/I4074/net049	net926	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4074/T4	vss	I0/I4074/net13	I0/I4074/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4074/T5	I0/I4074/net13	I0/I4074/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4074/T2	BL36	net926	I0/I4074/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4170/T3	I0/I4170/net049	net926	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4234/T5	I0/I4234/net13	I0/I4234/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4234/T2	BL39	net926	I0/I4234/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4202/T3	I0/I4202/net049	net926	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4202/T4	vss	I0/I4202/net13	I0/I4202/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4202/T5	I0/I4202/net13	I0/I4202/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4202/T2	BL38	net926	I0/I4202/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4169/T4	vss	I0/I4169/net13	I0/I4169/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4169/T5	I0/I4169/net13	I0/I4169/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4169/T2	BL37	net925	I0/I4169/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4073/T3	I0/I4073/net049	net925	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4073/T4	vss	I0/I4073/net13	I0/I4073/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4073/T5	I0/I4073/net13	I0/I4073/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4073/T2	BL36	net925	I0/I4073/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4169/T3	I0/I4169/net049	net925	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4233/T5	I0/I4233/net13	I0/I4233/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4233/T2	BL39	net925	I0/I4233/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4201/T3	I0/I4201/net049	net925	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4201/T4	vss	I0/I4201/net13	I0/I4201/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4201/T5	I0/I4201/net13	I0/I4201/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4201/T2	BL38	net925	I0/I4201/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4146/T4	vss	I0/I4146/net13	I0/I4146/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4146/T5	I0/I4146/net13	I0/I4146/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4146/T2	BL37	net924	I0/I4146/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4050/T3	I0/I4050/net049	net924	BL36bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4050/T4	vss	I0/I4050/net13	I0/I4050/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4050/T5	I0/I4050/net13	I0/I4050/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4050/T2	BL36	net924	I0/I4050/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4146/T3	I0/I4146/net049	net924	BL37bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4210/T5	I0/I4210/net13	I0/I4210/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4210/T2	BL39	net924	I0/I4210/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4178/T3	I0/I4178/net049	net924	BL38bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4178/T4	vss	I0/I4178/net13	I0/I4178/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4178/T5	I0/I4178/net13	I0/I4178/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4178/T2	BL38	net924	I0/I4178/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI109/T1	BL39	y4	p10	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI110/T1	p10bar	y3	BL38bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI111/T1	BL38	y3	p10	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI112/T1	p10bar	y2	BL37bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI113/T1	BL37	y2	p10	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI114/T1	p10bar	y1	BL36bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI115/T1	BL36	y1	p10	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T19	I32/net7	p9	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T18	p9bar	net680	I32/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T2	I11/net23	p10	I11/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T3	I11/net20	p10bar	I11/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T4	vss	vdd	I11/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T8	vss	I11/net20	I11/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T7	data9	I11/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T11	I33/net23	data9	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T16	I33/net15	net680	p10	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T17	vss	I33/net23	I33/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T19	I33/net7	p10	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T18	p10bar	net680	I33/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3932/T3	I0/I3932/net049	net955	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3932/T4	vss	I0/I3932/net13	I0/I3932/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3932/T5	I0/I3932/net13	I0/I3932/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3932/T2	BL32	net955	I0/I3932/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4220/T3	I0/I4220/net049	net955	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4220/T4	vss	I0/I4220/net13	I0/I4220/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3924/T3	I0/I3924/net049	net954	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3924/T4	vss	I0/I3924/net13	I0/I3924/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3924/T5	I0/I3924/net13	I0/I3924/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3924/T2	BL32	net954	I0/I3924/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4212/T3	I0/I4212/net049	net954	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4212/T4	vss	I0/I4212/net13	I0/I4212/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3923/T3	I0/I3923/net049	net953	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3923/T4	vss	I0/I3923/net13	I0/I3923/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3923/T5	I0/I3923/net13	I0/I3923/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3923/T2	BL32	net953	I0/I3923/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4211/T3	I0/I4211/net049	net953	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4211/T4	vss	I0/I4211/net13	I0/I4211/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3948/T3	I0/I3948/net049	net952	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3948/T4	vss	I0/I3948/net13	I0/I3948/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3948/T5	I0/I3948/net13	I0/I3948/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3948/T2	BL32	net952	I0/I3948/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4236/T3	I0/I4236/net049	net952	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4236/T4	vss	I0/I4236/net13	I0/I4236/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3929/T3	I0/I3929/net049	net951	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3929/T4	vss	I0/I3929/net13	I0/I3929/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3929/T5	I0/I3929/net13	I0/I3929/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3929/T2	BL32	net951	I0/I3929/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4217/T3	I0/I4217/net049	net951	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4217/T4	vss	I0/I4217/net13	I0/I4217/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3944/T3	I0/I3944/net049	net950	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3944/T4	vss	I0/I3944/net13	I0/I3944/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3944/T5	I0/I3944/net13	I0/I3944/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3944/T2	BL32	net950	I0/I3944/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4232/T3	I0/I4232/net049	net950	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4232/T4	vss	I0/I4232/net13	I0/I4232/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3942/T3	I0/I3942/net049	net949	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3942/T4	vss	I0/I3942/net13	I0/I3942/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3942/T5	I0/I3942/net13	I0/I3942/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3942/T2	BL32	net949	I0/I3942/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4230/T3	I0/I4230/net049	net949	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4230/T4	vss	I0/I4230/net13	I0/I4230/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3938/T3	I0/I3938/net049	net948	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3938/T4	vss	I0/I3938/net13	I0/I3938/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3938/T5	I0/I3938/net13	I0/I3938/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3938/T2	BL32	net948	I0/I3938/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4226/T3	I0/I4226/net049	net948	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4226/T4	vss	I0/I4226/net13	I0/I4226/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3930/T3	I0/I3930/net049	net947	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3930/T4	vss	I0/I3930/net13	I0/I3930/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3930/T5	I0/I3930/net13	I0/I3930/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3930/T2	BL32	net947	I0/I3930/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4218/T3	I0/I4218/net049	net947	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4218/T4	vss	I0/I4218/net13	I0/I4218/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3964/T2	BL33	net955	I0/I3964/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3956/T2	BL33	net954	I0/I3956/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3955/T2	BL33	net953	I0/I3955/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3980/T2	BL33	net952	I0/I3980/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3961/T2	BL33	net951	I0/I3961/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3976/T2	BL33	net950	I0/I3976/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3974/T2	BL33	net949	I0/I3974/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3970/T2	BL33	net948	I0/I3970/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3962/T2	BL33	net947	I0/I3962/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3964/T3	I0/I3964/net049	net955	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3956/T3	I0/I3956/net049	net954	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3964/T4	vss	I0/I3964/net13	I0/I3964/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3956/T4	vss	I0/I3956/net13	I0/I3956/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3964/T5	I0/I3964/net13	I0/I3964/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3956/T5	I0/I3956/net13	I0/I3956/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3955/T3	I0/I3955/net049	net953	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3980/T3	I0/I3980/net049	net952	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3955/T4	vss	I0/I3955/net13	I0/I3955/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3980/T4	vss	I0/I3980/net13	I0/I3980/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3955/T5	I0/I3955/net13	I0/I3955/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3980/T5	I0/I3980/net13	I0/I3980/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3961/T3	I0/I3961/net049	net951	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3961/T4	vss	I0/I3961/net13	I0/I3961/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3961/T5	I0/I3961/net13	I0/I3961/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3976/T3	I0/I3976/net049	net950	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3974/T3	I0/I3974/net049	net949	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3976/T4	vss	I0/I3976/net13	I0/I3976/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3974/T4	vss	I0/I3974/net13	I0/I3974/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3976/T5	I0/I3976/net13	I0/I3976/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3974/T5	I0/I3974/net13	I0/I3974/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3970/T3	I0/I3970/net049	net948	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3962/T3	I0/I3962/net049	net947	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3970/T4	vss	I0/I3970/net13	I0/I3970/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3962/T4	vss	I0/I3962/net13	I0/I3962/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3970/T5	I0/I3970/net13	I0/I3970/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3962/T5	I0/I3962/net13	I0/I3962/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3996/T2	BL34	net955	I0/I3996/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3988/T2	BL34	net954	I0/I3988/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3987/T2	BL34	net953	I0/I3987/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4012/T2	BL34	net952	I0/I4012/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3993/T2	BL34	net951	I0/I3993/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4008/T2	BL34	net950	I0/I4008/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4006/T2	BL34	net949	I0/I4006/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4002/T2	BL34	net948	I0/I4002/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3994/T2	BL34	net947	I0/I3994/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3996/T5	I0/I3996/net13	I0/I3996/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3988/T5	I0/I3988/net13	I0/I3988/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3987/T5	I0/I3987/net13	I0/I3987/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4012/T5	I0/I4012/net13	I0/I4012/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3993/T5	I0/I3993/net13	I0/I3993/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4008/T5	I0/I4008/net13	I0/I4008/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4006/T5	I0/I4006/net13	I0/I4006/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4002/T5	I0/I4002/net13	I0/I4002/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3994/T5	I0/I3994/net13	I0/I3994/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3996/T4	vss	I0/I3996/net13	I0/I3996/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3988/T4	vss	I0/I3988/net13	I0/I3988/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3987/T4	vss	I0/I3987/net13	I0/I3987/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4012/T4	vss	I0/I4012/net13	I0/I4012/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3993/T4	vss	I0/I3993/net13	I0/I3993/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4008/T4	vss	I0/I4008/net13	I0/I4008/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4006/T4	vss	I0/I4006/net13	I0/I4006/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4002/T4	vss	I0/I4002/net13	I0/I4002/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3994/T4	vss	I0/I3994/net13	I0/I3994/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3996/T3	I0/I3996/net049	net955	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3988/T3	I0/I3988/net049	net954	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3987/T3	I0/I3987/net049	net953	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4012/T3	I0/I4012/net049	net952	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3993/T3	I0/I3993/net049	net951	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4008/T3	I0/I4008/net049	net950	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4006/T3	I0/I4006/net049	net949	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4002/T3	I0/I4002/net049	net948	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3994/T3	I0/I3994/net049	net947	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3931/T3	I0/I3931/net049	net946	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3931/T4	vss	I0/I3931/net13	I0/I3931/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3931/T5	I0/I3931/net13	I0/I3931/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3931/T2	BL32	net946	I0/I3931/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4219/T3	I0/I4219/net049	net946	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4219/T4	vss	I0/I4219/net13	I0/I4219/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3921/T3	I0/I3921/net049	net945	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3921/T4	vss	I0/I3921/net13	I0/I3921/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3921/T5	I0/I3921/net13	I0/I3921/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3921/T2	BL32	net945	I0/I3921/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4209/T3	I0/I4209/net049	net945	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4209/T4	vss	I0/I4209/net13	I0/I4209/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3947/T3	I0/I3947/net049	net944	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3947/T4	vss	I0/I3947/net13	I0/I3947/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3947/T5	I0/I3947/net13	I0/I3947/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3947/T2	BL32	net944	I0/I3947/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4235/T3	I0/I4235/net049	net944	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4235/T4	vss	I0/I4235/net13	I0/I4235/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3941/T3	I0/I3941/net049	net943	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3941/T4	vss	I0/I3941/net13	I0/I3941/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3941/T5	I0/I3941/net13	I0/I3941/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3941/T2	BL32	net943	I0/I3941/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4229/T3	I0/I4229/net049	net943	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4229/T4	vss	I0/I4229/net13	I0/I4229/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3927/T3	I0/I3927/net049	net942	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3927/T4	vss	I0/I3927/net13	I0/I3927/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3927/T5	I0/I3927/net13	I0/I3927/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3927/T2	BL32	net942	I0/I3927/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4215/T3	I0/I4215/net049	net942	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4215/T4	vss	I0/I4215/net13	I0/I4215/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3920/T3	I0/I3920/net049	net941	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3920/T4	vss	I0/I3920/net13	I0/I3920/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3920/T5	I0/I3920/net13	I0/I3920/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3920/T2	BL32	net941	I0/I3920/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4208/T3	I0/I4208/net049	net941	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4208/T4	vss	I0/I4208/net13	I0/I4208/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3943/T3	I0/I3943/net049	net940	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3943/T4	vss	I0/I3943/net13	I0/I3943/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3943/T5	I0/I3943/net13	I0/I3943/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3943/T2	BL32	net940	I0/I3943/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4231/T3	I0/I4231/net049	net940	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4231/T4	vss	I0/I4231/net13	I0/I4231/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3940/T3	I0/I3940/net049	net939	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3940/T4	vss	I0/I3940/net13	I0/I3940/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3940/T5	I0/I3940/net13	I0/I3940/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3940/T2	BL32	net939	I0/I3940/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4228/T3	I0/I4228/net049	net939	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4228/T4	vss	I0/I4228/net13	I0/I4228/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3918/T3	I0/I3918/net049	net938	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3918/T4	vss	I0/I3918/net13	I0/I3918/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3918/T5	I0/I3918/net13	I0/I3918/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3918/T2	BL32	net938	I0/I3918/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4206/T3	I0/I4206/net049	net938	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4206/T4	vss	I0/I4206/net13	I0/I4206/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3963/T2	BL33	net946	I0/I3963/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3953/T2	BL33	net945	I0/I3953/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3979/T2	BL33	net944	I0/I3979/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3973/T2	BL33	net943	I0/I3973/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3959/T2	BL33	net942	I0/I3959/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3952/T2	BL33	net941	I0/I3952/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3975/T2	BL33	net940	I0/I3975/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3972/T2	BL33	net939	I0/I3972/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3950/T2	BL33	net938	I0/I3950/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3963/T3	I0/I3963/net049	net946	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3953/T3	I0/I3953/net049	net945	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3963/T4	vss	I0/I3963/net13	I0/I3963/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3953/T4	vss	I0/I3953/net13	I0/I3953/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3963/T5	I0/I3963/net13	I0/I3963/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3953/T5	I0/I3953/net13	I0/I3953/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3979/T3	I0/I3979/net049	net944	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3973/T3	I0/I3973/net049	net943	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3979/T4	vss	I0/I3979/net13	I0/I3979/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3973/T4	vss	I0/I3973/net13	I0/I3973/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3979/T5	I0/I3979/net13	I0/I3979/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3973/T5	I0/I3973/net13	I0/I3973/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3959/T3	I0/I3959/net049	net942	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3959/T4	vss	I0/I3959/net13	I0/I3959/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3959/T5	I0/I3959/net13	I0/I3959/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3952/T3	I0/I3952/net049	net941	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3975/T3	I0/I3975/net049	net940	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3952/T4	vss	I0/I3952/net13	I0/I3952/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3975/T4	vss	I0/I3975/net13	I0/I3975/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3952/T5	I0/I3952/net13	I0/I3952/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3975/T5	I0/I3975/net13	I0/I3975/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3972/T3	I0/I3972/net049	net939	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3950/T3	I0/I3950/net049	net938	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3972/T4	vss	I0/I3972/net13	I0/I3972/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3950/T4	vss	I0/I3950/net13	I0/I3950/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3972/T5	I0/I3972/net13	I0/I3972/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3950/T5	I0/I3950/net13	I0/I3950/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3995/T2	BL34	net946	I0/I3995/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3985/T2	BL34	net945	I0/I3985/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4011/T2	BL34	net944	I0/I4011/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4005/T2	BL34	net943	I0/I4005/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3991/T2	BL34	net942	I0/I3991/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3984/T2	BL34	net941	I0/I3984/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4007/T2	BL34	net940	I0/I4007/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4004/T2	BL34	net939	I0/I4004/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3982/T2	BL34	net938	I0/I3982/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3995/T5	I0/I3995/net13	I0/I3995/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3985/T5	I0/I3985/net13	I0/I3985/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4011/T5	I0/I4011/net13	I0/I4011/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4005/T5	I0/I4005/net13	I0/I4005/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3991/T5	I0/I3991/net13	I0/I3991/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3984/T5	I0/I3984/net13	I0/I3984/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4007/T5	I0/I4007/net13	I0/I4007/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4004/T5	I0/I4004/net13	I0/I4004/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3982/T5	I0/I3982/net13	I0/I3982/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3995/T4	vss	I0/I3995/net13	I0/I3995/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3985/T4	vss	I0/I3985/net13	I0/I3985/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4011/T4	vss	I0/I4011/net13	I0/I4011/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4005/T4	vss	I0/I4005/net13	I0/I4005/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3991/T4	vss	I0/I3991/net13	I0/I3991/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3984/T4	vss	I0/I3984/net13	I0/I3984/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4007/T4	vss	I0/I4007/net13	I0/I4007/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4004/T4	vss	I0/I4004/net13	I0/I4004/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3982/T4	vss	I0/I3982/net13	I0/I3982/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3995/T3	I0/I3995/net049	net946	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3985/T3	I0/I3985/net049	net945	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4011/T3	I0/I4011/net049	net944	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4005/T3	I0/I4005/net049	net943	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3991/T3	I0/I3991/net049	net942	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3984/T3	I0/I3984/net049	net941	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4007/T3	I0/I4007/net049	net940	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4004/T3	I0/I4004/net049	net939	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3982/T3	I0/I3982/net049	net938	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3919/T3	I0/I3919/net049	net937	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3919/T4	vss	I0/I3919/net13	I0/I3919/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3919/T5	I0/I3919/net13	I0/I3919/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3919/T2	BL32	net937	I0/I3919/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4207/T3	I0/I4207/net049	net937	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4207/T4	vss	I0/I4207/net13	I0/I4207/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3951/T2	BL33	net937	I0/I3951/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3983/T3	I0/I3983/net049	net937	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3983/T4	vss	I0/I3983/net13	I0/I3983/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3983/T5	I0/I3983/net13	I0/I3983/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3983/T2	BL34	net937	I0/I3983/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3951/T3	I0/I3951/net049	net937	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3951/T4	vss	I0/I3951/net13	I0/I3951/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3951/T5	I0/I3951/net13	I0/I3951/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3926/T3	I0/I3926/net049	net936	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3926/T4	vss	I0/I3926/net13	I0/I3926/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3926/T5	I0/I3926/net13	I0/I3926/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3926/T2	BL32	net936	I0/I3926/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4214/T3	I0/I4214/net049	net936	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4214/T4	vss	I0/I4214/net13	I0/I4214/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3958/T2	BL33	net936	I0/I3958/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3990/T3	I0/I3990/net049	net936	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3990/T4	vss	I0/I3990/net13	I0/I3990/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3990/T5	I0/I3990/net13	I0/I3990/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3990/T2	BL34	net936	I0/I3990/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3958/T3	I0/I3958/net049	net936	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3958/T4	vss	I0/I3958/net13	I0/I3958/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3958/T5	I0/I3958/net13	I0/I3958/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3928/T3	I0/I3928/net049	net935	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3928/T4	vss	I0/I3928/net13	I0/I3928/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3928/T5	I0/I3928/net13	I0/I3928/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3928/T2	BL32	net935	I0/I3928/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4216/T3	I0/I4216/net049	net935	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4216/T4	vss	I0/I4216/net13	I0/I4216/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3960/T2	BL33	net935	I0/I3960/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3992/T3	I0/I3992/net049	net935	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3992/T4	vss	I0/I3992/net13	I0/I3992/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3992/T5	I0/I3992/net13	I0/I3992/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3992/T2	BL34	net935	I0/I3992/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3960/T3	I0/I3960/net049	net935	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3960/T4	vss	I0/I3960/net13	I0/I3960/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3960/T5	I0/I3960/net13	I0/I3960/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3934/T3	I0/I3934/net049	net934	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3934/T4	vss	I0/I3934/net13	I0/I3934/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3934/T5	I0/I3934/net13	I0/I3934/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3934/T2	BL32	net934	I0/I3934/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4222/T3	I0/I4222/net049	net934	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4222/T4	vss	I0/I4222/net13	I0/I4222/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3966/T2	BL33	net934	I0/I3966/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3998/T3	I0/I3998/net049	net934	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3998/T4	vss	I0/I3998/net13	I0/I3998/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3998/T5	I0/I3998/net13	I0/I3998/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3998/T2	BL34	net934	I0/I3998/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3966/T3	I0/I3966/net049	net934	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3966/T4	vss	I0/I3966/net13	I0/I3966/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3966/T5	I0/I3966/net13	I0/I3966/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3936/T3	I0/I3936/net049	net933	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3936/T4	vss	I0/I3936/net13	I0/I3936/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3936/T5	I0/I3936/net13	I0/I3936/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3936/T2	BL32	net933	I0/I3936/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4224/T3	I0/I4224/net049	net933	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4224/T4	vss	I0/I4224/net13	I0/I4224/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3968/T2	BL33	net933	I0/I3968/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4000/T3	I0/I4000/net049	net933	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4000/T4	vss	I0/I4000/net13	I0/I4000/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4000/T5	I0/I4000/net13	I0/I4000/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4000/T2	BL34	net933	I0/I4000/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3968/T3	I0/I3968/net049	net933	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3968/T4	vss	I0/I3968/net13	I0/I3968/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3968/T5	I0/I3968/net13	I0/I3968/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3925/T3	I0/I3925/net049	net932	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3925/T4	vss	I0/I3925/net13	I0/I3925/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3925/T5	I0/I3925/net13	I0/I3925/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3925/T2	BL32	net932	I0/I3925/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4213/T3	I0/I4213/net049	net932	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4213/T4	vss	I0/I4213/net13	I0/I4213/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3957/T2	BL33	net932	I0/I3957/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3989/T3	I0/I3989/net049	net932	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3989/T4	vss	I0/I3989/net13	I0/I3989/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3989/T5	I0/I3989/net13	I0/I3989/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3989/T2	BL34	net932	I0/I3989/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3957/T3	I0/I3957/net049	net932	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3957/T4	vss	I0/I3957/net13	I0/I3957/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3957/T5	I0/I3957/net13	I0/I3957/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3939/T3	I0/I3939/net049	net931	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3939/T4	vss	I0/I3939/net13	I0/I3939/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3939/T5	I0/I3939/net13	I0/I3939/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3939/T2	BL32	net931	I0/I3939/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4227/T3	I0/I4227/net049	net931	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4227/T4	vss	I0/I4227/net13	I0/I4227/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3971/T2	BL33	net931	I0/I3971/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4003/T3	I0/I4003/net049	net931	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4003/T4	vss	I0/I4003/net13	I0/I4003/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4003/T5	I0/I4003/net13	I0/I4003/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4003/T2	BL34	net931	I0/I4003/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3971/T3	I0/I3971/net049	net931	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3971/T4	vss	I0/I3971/net13	I0/I3971/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3971/T5	I0/I3971/net13	I0/I3971/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3933/T3	I0/I3933/net049	net930	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3933/T4	vss	I0/I3933/net13	I0/I3933/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3933/T5	I0/I3933/net13	I0/I3933/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3933/T2	BL32	net930	I0/I3933/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4221/T3	I0/I4221/net049	net930	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4221/T4	vss	I0/I4221/net13	I0/I4221/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3965/T2	BL33	net930	I0/I3965/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3997/T3	I0/I3997/net049	net930	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3997/T4	vss	I0/I3997/net13	I0/I3997/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3997/T5	I0/I3997/net13	I0/I3997/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3997/T2	BL34	net930	I0/I3997/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3965/T3	I0/I3965/net049	net930	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3965/T4	vss	I0/I3965/net13	I0/I3965/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3965/T5	I0/I3965/net13	I0/I3965/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3937/T3	I0/I3937/net049	net929	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3937/T4	vss	I0/I3937/net13	I0/I3937/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3937/T5	I0/I3937/net13	I0/I3937/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3937/T2	BL32	net929	I0/I3937/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4225/T3	I0/I4225/net049	net929	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4225/T4	vss	I0/I4225/net13	I0/I4225/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3969/T2	BL33	net929	I0/I3969/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4001/T3	I0/I4001/net049	net929	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4001/T4	vss	I0/I4001/net13	I0/I4001/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4001/T5	I0/I4001/net13	I0/I4001/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4001/T2	BL34	net929	I0/I4001/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3969/T3	I0/I3969/net049	net929	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3969/T4	vss	I0/I3969/net13	I0/I3969/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3969/T5	I0/I3969/net13	I0/I3969/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3949/T3	I0/I3949/net049	net928	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3949/T4	vss	I0/I3949/net13	I0/I3949/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3949/T5	I0/I3949/net13	I0/I3949/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3949/T2	BL32	net928	I0/I3949/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4237/T3	I0/I4237/net049	net928	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4237/T4	vss	I0/I4237/net13	I0/I4237/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3981/T2	BL33	net928	I0/I3981/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4013/T3	I0/I4013/net049	net928	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4013/T4	vss	I0/I4013/net13	I0/I4013/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4013/T5	I0/I4013/net13	I0/I4013/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4013/T2	BL34	net928	I0/I4013/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3981/T3	I0/I3981/net049	net928	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3981/T4	vss	I0/I3981/net13	I0/I3981/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3981/T5	I0/I3981/net13	I0/I3981/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3935/T3	I0/I3935/net049	net927	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3935/T4	vss	I0/I3935/net13	I0/I3935/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3935/T5	I0/I3935/net13	I0/I3935/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3935/T2	BL32	net927	I0/I3935/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4223/T3	I0/I4223/net049	net927	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4223/T4	vss	I0/I4223/net13	I0/I4223/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3967/T2	BL33	net927	I0/I3967/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3999/T3	I0/I3999/net049	net927	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3999/T4	vss	I0/I3999/net13	I0/I3999/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3999/T5	I0/I3999/net13	I0/I3999/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3999/T2	BL34	net927	I0/I3999/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3967/T3	I0/I3967/net049	net927	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3967/T4	vss	I0/I3967/net13	I0/I3967/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3967/T5	I0/I3967/net13	I0/I3967/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3946/T3	I0/I3946/net049	net926	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3946/T4	vss	I0/I3946/net13	I0/I3946/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3946/T5	I0/I3946/net13	I0/I3946/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3946/T2	BL32	net926	I0/I3946/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4234/T3	I0/I4234/net049	net926	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4234/T4	vss	I0/I4234/net13	I0/I4234/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3978/T2	BL33	net926	I0/I3978/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4010/T3	I0/I4010/net049	net926	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4010/T4	vss	I0/I4010/net13	I0/I4010/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4010/T5	I0/I4010/net13	I0/I4010/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4010/T2	BL34	net926	I0/I4010/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3978/T3	I0/I3978/net049	net926	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3978/T4	vss	I0/I3978/net13	I0/I3978/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3978/T5	I0/I3978/net13	I0/I3978/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3945/T3	I0/I3945/net049	net925	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3945/T4	vss	I0/I3945/net13	I0/I3945/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3945/T5	I0/I3945/net13	I0/I3945/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3945/T2	BL32	net925	I0/I3945/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4233/T3	I0/I4233/net049	net925	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4233/T4	vss	I0/I4233/net13	I0/I4233/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3977/T2	BL33	net925	I0/I3977/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4009/T3	I0/I4009/net049	net925	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4009/T4	vss	I0/I4009/net13	I0/I4009/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4009/T5	I0/I4009/net13	I0/I4009/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4009/T2	BL34	net925	I0/I4009/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3977/T3	I0/I3977/net049	net925	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3977/T4	vss	I0/I3977/net13	I0/I3977/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3977/T5	I0/I3977/net13	I0/I3977/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3922/T3	I0/I3922/net049	net924	BL32bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3922/T4	vss	I0/I3922/net13	I0/I3922/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3922/T5	I0/I3922/net13	I0/I3922/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3922/T2	BL32	net924	I0/I3922/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4210/T3	I0/I4210/net049	net924	BL39bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4210/T4	vss	I0/I4210/net13	I0/I4210/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3954/T2	BL33	net924	I0/I3954/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3986/T3	I0/I3986/net049	net924	BL34bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3986/T4	vss	I0/I3986/net13	I0/I3986/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3986/T5	I0/I3986/net13	I0/I3986/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3986/T2	BL34	net924	I0/I3986/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3954/T3	I0/I3954/net049	net924	BL33bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3954/T4	vss	I0/I3954/net13	I0/I3954/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3954/T5	I0/I3954/net13	I0/I3954/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI102/T1	p9bar	y3	BL34bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI103/T1	BL34	y3	p9	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI104/T1	p9bar	y2	BL33bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI105/T1	BL33	y2	p9	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI106/T1	p9bar	y1	BL32bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI107/T1	BL32	y1	p9	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI108/T1	p10bar	y4	BL39bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T16	I31/net15	net680	p8	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T17	vss	I31/net23	I31/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T19	I31/net7	p8	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T18	p8bar	net680	I31/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T2	I10/net23	p9	I10/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T3	I10/net20	p9bar	I10/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T4	vss	vdd	I10/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T8	vss	I10/net20	I10/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T7	data8	I10/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T11	I32/net23	data8	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T16	I32/net15	net680	p9	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T17	vss	I32/net23	I32/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4028/T2	BL35	net955	I0/I4028/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4020/T2	BL35	net954	I0/I4020/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4019/T2	BL35	net953	I0/I4019/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4044/T2	BL35	net952	I0/I4044/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4025/T2	BL35	net951	I0/I4025/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4040/T2	BL35	net950	I0/I4040/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4038/T2	BL35	net949	I0/I4038/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4034/T2	BL35	net948	I0/I4034/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4026/T2	BL35	net947	I0/I4026/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4028/T5	I0/I4028/net13	I0/I4028/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4020/T5	I0/I4020/net13	I0/I4020/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4019/T5	I0/I4019/net13	I0/I4019/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4044/T5	I0/I4044/net13	I0/I4044/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4025/T5	I0/I4025/net13	I0/I4025/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4040/T5	I0/I4040/net13	I0/I4040/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4038/T5	I0/I4038/net13	I0/I4038/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4034/T5	I0/I4034/net13	I0/I4034/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4026/T5	I0/I4026/net13	I0/I4026/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4028/T4	vss	I0/I4028/net13	I0/I4028/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4020/T4	vss	I0/I4020/net13	I0/I4020/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4019/T4	vss	I0/I4019/net13	I0/I4019/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4044/T4	vss	I0/I4044/net13	I0/I4044/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4025/T4	vss	I0/I4025/net13	I0/I4025/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4040/T4	vss	I0/I4040/net13	I0/I4040/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4038/T4	vss	I0/I4038/net13	I0/I4038/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4034/T4	vss	I0/I4034/net13	I0/I4034/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4026/T4	vss	I0/I4026/net13	I0/I4026/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4028/T3	I0/I4028/net049	net955	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4020/T3	I0/I4020/net049	net954	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4019/T3	I0/I4019/net049	net953	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4044/T3	I0/I4044/net049	net952	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4025/T3	I0/I4025/net049	net951	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4040/T3	I0/I4040/net049	net950	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4038/T3	I0/I4038/net049	net949	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4034/T3	I0/I4034/net049	net948	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4026/T3	I0/I4026/net049	net947	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3804/T4	vss	I0/I3804/net13	I0/I3804/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3796/T4	vss	I0/I3796/net13	I0/I3796/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3804/T5	I0/I3804/net13	I0/I3804/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3796/T5	I0/I3796/net13	I0/I3796/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3804/T2	BL28	net955	I0/I3804/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3796/T2	BL28	net954	I0/I3796/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3795/T4	vss	I0/I3795/net13	I0/I3795/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3820/T4	vss	I0/I3820/net13	I0/I3820/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3795/T5	I0/I3795/net13	I0/I3795/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3820/T5	I0/I3820/net13	I0/I3820/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3795/T2	BL28	net953	I0/I3795/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3820/T2	BL28	net952	I0/I3820/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3801/T4	vss	I0/I3801/net13	I0/I3801/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3801/T5	I0/I3801/net13	I0/I3801/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3801/T2	BL28	net951	I0/I3801/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3816/T4	vss	I0/I3816/net13	I0/I3816/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3814/T4	vss	I0/I3814/net13	I0/I3814/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3816/T5	I0/I3816/net13	I0/I3816/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3814/T5	I0/I3814/net13	I0/I3814/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3816/T2	BL28	net950	I0/I3816/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3814/T2	BL28	net949	I0/I3814/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3810/T4	vss	I0/I3810/net13	I0/I3810/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3802/T4	vss	I0/I3802/net13	I0/I3802/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3810/T5	I0/I3810/net13	I0/I3810/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3802/T5	I0/I3802/net13	I0/I3802/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3810/T2	BL28	net948	I0/I3810/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3802/T2	BL28	net947	I0/I3802/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3804/T3	I0/I3804/net049	net955	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3796/T3	I0/I3796/net049	net954	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3795/T3	I0/I3795/net049	net953	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3820/T3	I0/I3820/net049	net952	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3801/T3	I0/I3801/net049	net951	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3816/T3	I0/I3816/net049	net950	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3814/T3	I0/I3814/net049	net949	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3810/T3	I0/I3810/net049	net948	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3802/T3	I0/I3802/net049	net947	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3868/T5	I0/I3868/net13	I0/I3868/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3868/T2	BL30	net955	I0/I3868/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3836/T3	I0/I3836/net049	net955	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3836/T4	vss	I0/I3836/net13	I0/I3836/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3836/T5	I0/I3836/net13	I0/I3836/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3836/T2	BL29	net955	I0/I3836/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3860/T5	I0/I3860/net13	I0/I3860/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3860/T2	BL30	net954	I0/I3860/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3828/T3	I0/I3828/net049	net954	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3828/T4	vss	I0/I3828/net13	I0/I3828/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3828/T5	I0/I3828/net13	I0/I3828/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3828/T2	BL29	net954	I0/I3828/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3859/T5	I0/I3859/net13	I0/I3859/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3859/T2	BL30	net953	I0/I3859/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3827/T3	I0/I3827/net049	net953	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3827/T4	vss	I0/I3827/net13	I0/I3827/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3827/T5	I0/I3827/net13	I0/I3827/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3827/T2	BL29	net953	I0/I3827/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3884/T5	I0/I3884/net13	I0/I3884/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3884/T2	BL30	net952	I0/I3884/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3852/T3	I0/I3852/net049	net952	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3852/T4	vss	I0/I3852/net13	I0/I3852/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3852/T5	I0/I3852/net13	I0/I3852/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3852/T2	BL29	net952	I0/I3852/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3865/T5	I0/I3865/net13	I0/I3865/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3865/T2	BL30	net951	I0/I3865/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3833/T3	I0/I3833/net049	net951	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3833/T4	vss	I0/I3833/net13	I0/I3833/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3833/T5	I0/I3833/net13	I0/I3833/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3833/T2	BL29	net951	I0/I3833/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3880/T5	I0/I3880/net13	I0/I3880/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3880/T2	BL30	net950	I0/I3880/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3848/T3	I0/I3848/net049	net950	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3848/T4	vss	I0/I3848/net13	I0/I3848/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3848/T5	I0/I3848/net13	I0/I3848/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3848/T2	BL29	net950	I0/I3848/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3878/T5	I0/I3878/net13	I0/I3878/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3878/T2	BL30	net949	I0/I3878/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3846/T3	I0/I3846/net049	net949	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3846/T4	vss	I0/I3846/net13	I0/I3846/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3846/T5	I0/I3846/net13	I0/I3846/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3846/T2	BL29	net949	I0/I3846/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3874/T5	I0/I3874/net13	I0/I3874/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3874/T2	BL30	net948	I0/I3874/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3842/T3	I0/I3842/net049	net948	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3842/T4	vss	I0/I3842/net13	I0/I3842/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3842/T5	I0/I3842/net13	I0/I3842/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3842/T2	BL29	net948	I0/I3842/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3866/T5	I0/I3866/net13	I0/I3866/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3866/T2	BL30	net947	I0/I3866/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3834/T3	I0/I3834/net049	net947	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3834/T4	vss	I0/I3834/net13	I0/I3834/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3834/T5	I0/I3834/net13	I0/I3834/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3834/T2	BL29	net947	I0/I3834/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4027/T2	BL35	net946	I0/I4027/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4017/T2	BL35	net945	I0/I4017/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4043/T2	BL35	net944	I0/I4043/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4037/T2	BL35	net943	I0/I4037/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4023/T2	BL35	net942	I0/I4023/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4016/T2	BL35	net941	I0/I4016/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4039/T2	BL35	net940	I0/I4039/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4036/T2	BL35	net939	I0/I4036/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4014/T2	BL35	net938	I0/I4014/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4027/T5	I0/I4027/net13	I0/I4027/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4017/T5	I0/I4017/net13	I0/I4017/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4043/T5	I0/I4043/net13	I0/I4043/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4037/T5	I0/I4037/net13	I0/I4037/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4023/T5	I0/I4023/net13	I0/I4023/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4016/T5	I0/I4016/net13	I0/I4016/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4039/T5	I0/I4039/net13	I0/I4039/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4036/T5	I0/I4036/net13	I0/I4036/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4014/T5	I0/I4014/net13	I0/I4014/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4027/T4	vss	I0/I4027/net13	I0/I4027/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4017/T4	vss	I0/I4017/net13	I0/I4017/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4043/T4	vss	I0/I4043/net13	I0/I4043/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4037/T4	vss	I0/I4037/net13	I0/I4037/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4023/T4	vss	I0/I4023/net13	I0/I4023/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4016/T4	vss	I0/I4016/net13	I0/I4016/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4039/T4	vss	I0/I4039/net13	I0/I4039/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4036/T4	vss	I0/I4036/net13	I0/I4036/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4014/T4	vss	I0/I4014/net13	I0/I4014/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4027/T3	I0/I4027/net049	net946	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4017/T3	I0/I4017/net049	net945	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4043/T3	I0/I4043/net049	net944	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4037/T3	I0/I4037/net049	net943	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4023/T3	I0/I4023/net049	net942	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4016/T3	I0/I4016/net049	net941	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4039/T3	I0/I4039/net049	net940	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4036/T3	I0/I4036/net049	net939	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4014/T3	I0/I4014/net049	net938	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3803/T4	vss	I0/I3803/net13	I0/I3803/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3793/T4	vss	I0/I3793/net13	I0/I3793/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3803/T5	I0/I3803/net13	I0/I3803/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3793/T5	I0/I3793/net13	I0/I3793/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3803/T2	BL28	net946	I0/I3803/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3793/T2	BL28	net945	I0/I3793/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3819/T4	vss	I0/I3819/net13	I0/I3819/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3813/T4	vss	I0/I3813/net13	I0/I3813/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3819/T5	I0/I3819/net13	I0/I3819/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3813/T5	I0/I3813/net13	I0/I3813/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3819/T2	BL28	net944	I0/I3819/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3813/T2	BL28	net943	I0/I3813/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3799/T4	vss	I0/I3799/net13	I0/I3799/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3799/T5	I0/I3799/net13	I0/I3799/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3799/T2	BL28	net942	I0/I3799/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3792/T4	vss	I0/I3792/net13	I0/I3792/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3815/T4	vss	I0/I3815/net13	I0/I3815/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3792/T5	I0/I3792/net13	I0/I3792/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3815/T5	I0/I3815/net13	I0/I3815/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3792/T2	BL28	net941	I0/I3792/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3815/T2	BL28	net940	I0/I3815/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3812/T4	vss	I0/I3812/net13	I0/I3812/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3790/T4	vss	I0/I3790/net13	I0/I3790/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3812/T5	I0/I3812/net13	I0/I3812/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3790/T5	I0/I3790/net13	I0/I3790/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3812/T2	BL28	net939	I0/I3812/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3790/T2	BL28	net938	I0/I3790/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3803/T3	I0/I3803/net049	net946	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3793/T3	I0/I3793/net049	net945	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3819/T3	I0/I3819/net049	net944	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3813/T3	I0/I3813/net049	net943	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3799/T3	I0/I3799/net049	net942	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3792/T3	I0/I3792/net049	net941	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3815/T3	I0/I3815/net049	net940	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3812/T3	I0/I3812/net049	net939	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3790/T3	I0/I3790/net049	net938	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3867/T5	I0/I3867/net13	I0/I3867/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3867/T2	BL30	net946	I0/I3867/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3835/T3	I0/I3835/net049	net946	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3835/T4	vss	I0/I3835/net13	I0/I3835/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3835/T5	I0/I3835/net13	I0/I3835/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3835/T2	BL29	net946	I0/I3835/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3857/T5	I0/I3857/net13	I0/I3857/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3857/T2	BL30	net945	I0/I3857/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3825/T3	I0/I3825/net049	net945	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3825/T4	vss	I0/I3825/net13	I0/I3825/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3825/T5	I0/I3825/net13	I0/I3825/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3825/T2	BL29	net945	I0/I3825/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3883/T5	I0/I3883/net13	I0/I3883/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3883/T2	BL30	net944	I0/I3883/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3851/T3	I0/I3851/net049	net944	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3851/T4	vss	I0/I3851/net13	I0/I3851/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3851/T5	I0/I3851/net13	I0/I3851/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3851/T2	BL29	net944	I0/I3851/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3877/T5	I0/I3877/net13	I0/I3877/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3877/T2	BL30	net943	I0/I3877/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3845/T3	I0/I3845/net049	net943	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3845/T4	vss	I0/I3845/net13	I0/I3845/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3845/T5	I0/I3845/net13	I0/I3845/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3845/T2	BL29	net943	I0/I3845/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3863/T5	I0/I3863/net13	I0/I3863/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3863/T2	BL30	net942	I0/I3863/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3831/T3	I0/I3831/net049	net942	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3831/T4	vss	I0/I3831/net13	I0/I3831/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3831/T5	I0/I3831/net13	I0/I3831/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3831/T2	BL29	net942	I0/I3831/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3856/T5	I0/I3856/net13	I0/I3856/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3856/T2	BL30	net941	I0/I3856/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3824/T3	I0/I3824/net049	net941	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3824/T4	vss	I0/I3824/net13	I0/I3824/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3824/T5	I0/I3824/net13	I0/I3824/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3824/T2	BL29	net941	I0/I3824/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3879/T5	I0/I3879/net13	I0/I3879/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3879/T2	BL30	net940	I0/I3879/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3847/T3	I0/I3847/net049	net940	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3847/T4	vss	I0/I3847/net13	I0/I3847/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3847/T5	I0/I3847/net13	I0/I3847/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3847/T2	BL29	net940	I0/I3847/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3876/T5	I0/I3876/net13	I0/I3876/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3876/T2	BL30	net939	I0/I3876/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3844/T3	I0/I3844/net049	net939	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3844/T4	vss	I0/I3844/net13	I0/I3844/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3844/T5	I0/I3844/net13	I0/I3844/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3844/T2	BL29	net939	I0/I3844/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3854/T5	I0/I3854/net13	I0/I3854/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3854/T2	BL30	net938	I0/I3854/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3822/T3	I0/I3822/net049	net938	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3822/T4	vss	I0/I3822/net13	I0/I3822/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3822/T5	I0/I3822/net13	I0/I3822/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3822/T2	BL29	net938	I0/I3822/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3791/T4	vss	I0/I3791/net13	I0/I3791/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3791/T5	I0/I3791/net13	I0/I3791/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3791/T2	BL28	net937	I0/I3791/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4015/T3	I0/I4015/net049	net937	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4015/T4	vss	I0/I4015/net13	I0/I4015/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4015/T5	I0/I4015/net13	I0/I4015/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4015/T2	BL35	net937	I0/I4015/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3791/T3	I0/I3791/net049	net937	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3855/T5	I0/I3855/net13	I0/I3855/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3855/T2	BL30	net937	I0/I3855/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3823/T3	I0/I3823/net049	net937	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3823/T4	vss	I0/I3823/net13	I0/I3823/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3823/T5	I0/I3823/net13	I0/I3823/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3823/T2	BL29	net937	I0/I3823/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3798/T4	vss	I0/I3798/net13	I0/I3798/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3798/T5	I0/I3798/net13	I0/I3798/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3798/T2	BL28	net936	I0/I3798/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4022/T3	I0/I4022/net049	net936	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4022/T4	vss	I0/I4022/net13	I0/I4022/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4022/T5	I0/I4022/net13	I0/I4022/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4022/T2	BL35	net936	I0/I4022/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3798/T3	I0/I3798/net049	net936	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3862/T5	I0/I3862/net13	I0/I3862/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3862/T2	BL30	net936	I0/I3862/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3830/T3	I0/I3830/net049	net936	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3830/T4	vss	I0/I3830/net13	I0/I3830/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3830/T5	I0/I3830/net13	I0/I3830/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3830/T2	BL29	net936	I0/I3830/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3800/T4	vss	I0/I3800/net13	I0/I3800/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3800/T5	I0/I3800/net13	I0/I3800/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3800/T2	BL28	net935	I0/I3800/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4024/T3	I0/I4024/net049	net935	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4024/T4	vss	I0/I4024/net13	I0/I4024/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4024/T5	I0/I4024/net13	I0/I4024/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4024/T2	BL35	net935	I0/I4024/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3800/T3	I0/I3800/net049	net935	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3864/T5	I0/I3864/net13	I0/I3864/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3864/T2	BL30	net935	I0/I3864/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3832/T3	I0/I3832/net049	net935	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3832/T4	vss	I0/I3832/net13	I0/I3832/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3832/T5	I0/I3832/net13	I0/I3832/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3832/T2	BL29	net935	I0/I3832/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3806/T4	vss	I0/I3806/net13	I0/I3806/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3806/T5	I0/I3806/net13	I0/I3806/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3806/T2	BL28	net934	I0/I3806/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4030/T3	I0/I4030/net049	net934	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4030/T4	vss	I0/I4030/net13	I0/I4030/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4030/T5	I0/I4030/net13	I0/I4030/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4030/T2	BL35	net934	I0/I4030/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3806/T3	I0/I3806/net049	net934	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3870/T5	I0/I3870/net13	I0/I3870/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3870/T2	BL30	net934	I0/I3870/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3838/T3	I0/I3838/net049	net934	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3838/T4	vss	I0/I3838/net13	I0/I3838/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3838/T5	I0/I3838/net13	I0/I3838/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3838/T2	BL29	net934	I0/I3838/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3808/T4	vss	I0/I3808/net13	I0/I3808/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3808/T5	I0/I3808/net13	I0/I3808/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3808/T2	BL28	net933	I0/I3808/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4032/T3	I0/I4032/net049	net933	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4032/T4	vss	I0/I4032/net13	I0/I4032/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4032/T5	I0/I4032/net13	I0/I4032/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4032/T2	BL35	net933	I0/I4032/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3808/T3	I0/I3808/net049	net933	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3872/T5	I0/I3872/net13	I0/I3872/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3872/T2	BL30	net933	I0/I3872/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3840/T3	I0/I3840/net049	net933	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3840/T4	vss	I0/I3840/net13	I0/I3840/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3840/T5	I0/I3840/net13	I0/I3840/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3840/T2	BL29	net933	I0/I3840/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3797/T4	vss	I0/I3797/net13	I0/I3797/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3797/T5	I0/I3797/net13	I0/I3797/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3797/T2	BL28	net932	I0/I3797/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4021/T3	I0/I4021/net049	net932	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4021/T4	vss	I0/I4021/net13	I0/I4021/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4021/T5	I0/I4021/net13	I0/I4021/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4021/T2	BL35	net932	I0/I4021/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3797/T3	I0/I3797/net049	net932	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3861/T5	I0/I3861/net13	I0/I3861/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3861/T2	BL30	net932	I0/I3861/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3829/T3	I0/I3829/net049	net932	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3829/T4	vss	I0/I3829/net13	I0/I3829/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3829/T5	I0/I3829/net13	I0/I3829/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3829/T2	BL29	net932	I0/I3829/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3811/T4	vss	I0/I3811/net13	I0/I3811/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3811/T5	I0/I3811/net13	I0/I3811/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3811/T2	BL28	net931	I0/I3811/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4035/T3	I0/I4035/net049	net931	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4035/T4	vss	I0/I4035/net13	I0/I4035/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4035/T5	I0/I4035/net13	I0/I4035/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4035/T2	BL35	net931	I0/I4035/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3811/T3	I0/I3811/net049	net931	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3875/T5	I0/I3875/net13	I0/I3875/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3875/T2	BL30	net931	I0/I3875/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3843/T3	I0/I3843/net049	net931	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3843/T4	vss	I0/I3843/net13	I0/I3843/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3843/T5	I0/I3843/net13	I0/I3843/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3843/T2	BL29	net931	I0/I3843/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3805/T4	vss	I0/I3805/net13	I0/I3805/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3805/T5	I0/I3805/net13	I0/I3805/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3805/T2	BL28	net930	I0/I3805/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4029/T3	I0/I4029/net049	net930	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4029/T4	vss	I0/I4029/net13	I0/I4029/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4029/T5	I0/I4029/net13	I0/I4029/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4029/T2	BL35	net930	I0/I4029/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3805/T3	I0/I3805/net049	net930	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3869/T5	I0/I3869/net13	I0/I3869/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3869/T2	BL30	net930	I0/I3869/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3837/T3	I0/I3837/net049	net930	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3837/T4	vss	I0/I3837/net13	I0/I3837/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3837/T5	I0/I3837/net13	I0/I3837/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3837/T2	BL29	net930	I0/I3837/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3809/T4	vss	I0/I3809/net13	I0/I3809/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3809/T5	I0/I3809/net13	I0/I3809/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3809/T2	BL28	net929	I0/I3809/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4033/T3	I0/I4033/net049	net929	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4033/T4	vss	I0/I4033/net13	I0/I4033/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4033/T5	I0/I4033/net13	I0/I4033/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4033/T2	BL35	net929	I0/I4033/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3809/T3	I0/I3809/net049	net929	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3873/T5	I0/I3873/net13	I0/I3873/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3873/T2	BL30	net929	I0/I3873/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3841/T3	I0/I3841/net049	net929	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3841/T4	vss	I0/I3841/net13	I0/I3841/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3841/T5	I0/I3841/net13	I0/I3841/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3841/T2	BL29	net929	I0/I3841/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3821/T4	vss	I0/I3821/net13	I0/I3821/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3821/T5	I0/I3821/net13	I0/I3821/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3821/T2	BL28	net928	I0/I3821/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4045/T3	I0/I4045/net049	net928	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4045/T4	vss	I0/I4045/net13	I0/I4045/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4045/T5	I0/I4045/net13	I0/I4045/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4045/T2	BL35	net928	I0/I4045/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3821/T3	I0/I3821/net049	net928	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3885/T5	I0/I3885/net13	I0/I3885/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3885/T2	BL30	net928	I0/I3885/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3853/T3	I0/I3853/net049	net928	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3853/T4	vss	I0/I3853/net13	I0/I3853/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3853/T5	I0/I3853/net13	I0/I3853/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3853/T2	BL29	net928	I0/I3853/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3807/T4	vss	I0/I3807/net13	I0/I3807/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3807/T5	I0/I3807/net13	I0/I3807/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3807/T2	BL28	net927	I0/I3807/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4031/T3	I0/I4031/net049	net927	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4031/T4	vss	I0/I4031/net13	I0/I4031/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4031/T5	I0/I4031/net13	I0/I4031/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4031/T2	BL35	net927	I0/I4031/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3807/T3	I0/I3807/net049	net927	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3871/T5	I0/I3871/net13	I0/I3871/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3871/T2	BL30	net927	I0/I3871/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3839/T3	I0/I3839/net049	net927	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3839/T4	vss	I0/I3839/net13	I0/I3839/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3839/T5	I0/I3839/net13	I0/I3839/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3839/T2	BL29	net927	I0/I3839/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3818/T4	vss	I0/I3818/net13	I0/I3818/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3818/T5	I0/I3818/net13	I0/I3818/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3818/T2	BL28	net926	I0/I3818/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4042/T3	I0/I4042/net049	net926	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4042/T4	vss	I0/I4042/net13	I0/I4042/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4042/T5	I0/I4042/net13	I0/I4042/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4042/T2	BL35	net926	I0/I4042/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3818/T3	I0/I3818/net049	net926	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3882/T5	I0/I3882/net13	I0/I3882/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3882/T2	BL30	net926	I0/I3882/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3850/T3	I0/I3850/net049	net926	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3850/T4	vss	I0/I3850/net13	I0/I3850/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3850/T5	I0/I3850/net13	I0/I3850/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3850/T2	BL29	net926	I0/I3850/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3817/T4	vss	I0/I3817/net13	I0/I3817/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3817/T5	I0/I3817/net13	I0/I3817/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3817/T2	BL28	net925	I0/I3817/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4041/T3	I0/I4041/net049	net925	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4041/T4	vss	I0/I4041/net13	I0/I4041/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4041/T5	I0/I4041/net13	I0/I4041/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4041/T2	BL35	net925	I0/I4041/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3817/T3	I0/I3817/net049	net925	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3881/T5	I0/I3881/net13	I0/I3881/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3881/T2	BL30	net925	I0/I3881/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3849/T3	I0/I3849/net049	net925	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3849/T4	vss	I0/I3849/net13	I0/I3849/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3849/T5	I0/I3849/net13	I0/I3849/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3849/T2	BL29	net925	I0/I3849/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3794/T4	vss	I0/I3794/net13	I0/I3794/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3794/T5	I0/I3794/net13	I0/I3794/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3794/T2	BL28	net924	I0/I3794/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4018/T3	I0/I4018/net049	net924	BL35bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4018/T4	vss	I0/I4018/net13	I0/I4018/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4018/T5	I0/I4018/net13	I0/I4018/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4018/T2	BL35	net924	I0/I4018/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3794/T3	I0/I3794/net049	net924	BL28bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3858/T5	I0/I3858/net13	I0/I3858/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3858/T2	BL30	net924	I0/I3858/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3826/T3	I0/I3826/net049	net924	BL29bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3826/T4	vss	I0/I3826/net13	I0/I3826/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3826/T5	I0/I3826/net13	I0/I3826/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3826/T2	BL29	net924	I0/I3826/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T3	I8/net20	p8bar	I8/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T4	vss	vdd	I8/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI99/T1	BL28	y1	p8	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T8	vss	I8/net20	I8/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI100/T1	p9bar	y4	BL35bar	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T7	data7	I8/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T11	I31/net23	data7	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI101/T1	BL35	y4	p9	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T11	I29/net23	data6	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI95/T1	BL30	y3	p8	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T16	I29/net15	net680	p7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI96/T1	p8bar	y2	BL29bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T17	vss	I29/net23	I29/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T19	I29/net7	p7	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T18	p7bar	net680	I29/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI97/T1	BL29	y2	p8	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI98/T1	p8bar	y1	BL28bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T2	I8/net23	p8	I8/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3900/T3	I0/I3900/net049	net955	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3900/T4	vss	I0/I3900/net13	I0/I3900/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3900/T5	I0/I3900/net13	I0/I3900/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3900/T2	BL31	net955	I0/I3900/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3868/T3	I0/I3868/net049	net955	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3868/T4	vss	I0/I3868/net13	I0/I3868/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3892/T3	I0/I3892/net049	net954	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3892/T4	vss	I0/I3892/net13	I0/I3892/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3892/T5	I0/I3892/net13	I0/I3892/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3892/T2	BL31	net954	I0/I3892/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3860/T3	I0/I3860/net049	net954	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3860/T4	vss	I0/I3860/net13	I0/I3860/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3891/T3	I0/I3891/net049	net953	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3891/T4	vss	I0/I3891/net13	I0/I3891/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3891/T5	I0/I3891/net13	I0/I3891/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3891/T2	BL31	net953	I0/I3891/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3859/T3	I0/I3859/net049	net953	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3859/T4	vss	I0/I3859/net13	I0/I3859/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3916/T3	I0/I3916/net049	net952	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3916/T4	vss	I0/I3916/net13	I0/I3916/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3916/T5	I0/I3916/net13	I0/I3916/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3916/T2	BL31	net952	I0/I3916/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3884/T3	I0/I3884/net049	net952	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3884/T4	vss	I0/I3884/net13	I0/I3884/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3897/T3	I0/I3897/net049	net951	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3897/T4	vss	I0/I3897/net13	I0/I3897/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3897/T5	I0/I3897/net13	I0/I3897/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3897/T2	BL31	net951	I0/I3897/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3865/T3	I0/I3865/net049	net951	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3865/T4	vss	I0/I3865/net13	I0/I3865/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3912/T3	I0/I3912/net049	net950	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3912/T4	vss	I0/I3912/net13	I0/I3912/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3912/T5	I0/I3912/net13	I0/I3912/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3912/T2	BL31	net950	I0/I3912/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3880/T3	I0/I3880/net049	net950	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3880/T4	vss	I0/I3880/net13	I0/I3880/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3910/T3	I0/I3910/net049	net949	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3910/T4	vss	I0/I3910/net13	I0/I3910/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3910/T5	I0/I3910/net13	I0/I3910/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3910/T2	BL31	net949	I0/I3910/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3878/T3	I0/I3878/net049	net949	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3878/T4	vss	I0/I3878/net13	I0/I3878/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3906/T3	I0/I3906/net049	net948	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3906/T4	vss	I0/I3906/net13	I0/I3906/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3906/T5	I0/I3906/net13	I0/I3906/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3906/T2	BL31	net948	I0/I3906/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3874/T3	I0/I3874/net049	net948	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3874/T4	vss	I0/I3874/net13	I0/I3874/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3898/T3	I0/I3898/net049	net947	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3898/T4	vss	I0/I3898/net13	I0/I3898/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3898/T5	I0/I3898/net13	I0/I3898/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3898/T2	BL31	net947	I0/I3898/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3866/T3	I0/I3866/net049	net947	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3866/T4	vss	I0/I3866/net13	I0/I3866/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3676/T2	BL24	net955	I0/I3676/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3668/T2	BL24	net954	I0/I3668/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3667/T2	BL24	net953	I0/I3667/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3692/T2	BL24	net952	I0/I3692/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3673/T2	BL24	net951	I0/I3673/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3688/T2	BL24	net950	I0/I3688/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3686/T2	BL24	net949	I0/I3686/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3682/T2	BL24	net948	I0/I3682/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3674/T2	BL24	net947	I0/I3674/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3676/T3	I0/I3676/net049	net955	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3668/T3	I0/I3668/net049	net954	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3676/T4	vss	I0/I3676/net13	I0/I3676/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3668/T4	vss	I0/I3668/net13	I0/I3668/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3676/T5	I0/I3676/net13	I0/I3676/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3668/T5	I0/I3668/net13	I0/I3668/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3667/T3	I0/I3667/net049	net953	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3692/T3	I0/I3692/net049	net952	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3667/T4	vss	I0/I3667/net13	I0/I3667/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3692/T4	vss	I0/I3692/net13	I0/I3692/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3667/T5	I0/I3667/net13	I0/I3667/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3692/T5	I0/I3692/net13	I0/I3692/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3673/T3	I0/I3673/net049	net951	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3673/T4	vss	I0/I3673/net13	I0/I3673/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3673/T5	I0/I3673/net13	I0/I3673/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3688/T3	I0/I3688/net049	net950	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3686/T3	I0/I3686/net049	net949	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3688/T4	vss	I0/I3688/net13	I0/I3688/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3686/T4	vss	I0/I3686/net13	I0/I3686/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3688/T5	I0/I3688/net13	I0/I3688/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3686/T5	I0/I3686/net13	I0/I3686/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3682/T3	I0/I3682/net049	net948	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3674/T3	I0/I3674/net049	net947	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3682/T4	vss	I0/I3682/net13	I0/I3682/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3674/T4	vss	I0/I3674/net13	I0/I3674/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3682/T5	I0/I3682/net13	I0/I3682/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3674/T5	I0/I3674/net13	I0/I3674/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3708/T2	BL25	net955	I0/I3708/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3700/T2	BL25	net954	I0/I3700/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3699/T2	BL25	net953	I0/I3699/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3724/T2	BL25	net952	I0/I3724/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3705/T2	BL25	net951	I0/I3705/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3720/T2	BL25	net950	I0/I3720/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3718/T2	BL25	net949	I0/I3718/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3714/T2	BL25	net948	I0/I3714/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3706/T2	BL25	net947	I0/I3706/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3708/T5	I0/I3708/net13	I0/I3708/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3700/T5	I0/I3700/net13	I0/I3700/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3699/T5	I0/I3699/net13	I0/I3699/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3724/T5	I0/I3724/net13	I0/I3724/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3705/T5	I0/I3705/net13	I0/I3705/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3720/T5	I0/I3720/net13	I0/I3720/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3718/T5	I0/I3718/net13	I0/I3718/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3714/T5	I0/I3714/net13	I0/I3714/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3706/T5	I0/I3706/net13	I0/I3706/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3708/T4	vss	I0/I3708/net13	I0/I3708/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3700/T4	vss	I0/I3700/net13	I0/I3700/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3699/T4	vss	I0/I3699/net13	I0/I3699/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3724/T4	vss	I0/I3724/net13	I0/I3724/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3705/T4	vss	I0/I3705/net13	I0/I3705/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3720/T4	vss	I0/I3720/net13	I0/I3720/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3718/T4	vss	I0/I3718/net13	I0/I3718/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3714/T4	vss	I0/I3714/net13	I0/I3714/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3706/T4	vss	I0/I3706/net13	I0/I3706/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3708/T3	I0/I3708/net049	net955	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3700/T3	I0/I3700/net049	net954	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3699/T3	I0/I3699/net049	net953	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3724/T3	I0/I3724/net049	net952	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3705/T3	I0/I3705/net049	net951	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3720/T3	I0/I3720/net049	net950	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3718/T3	I0/I3718/net049	net949	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3714/T3	I0/I3714/net049	net948	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3706/T3	I0/I3706/net049	net947	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3899/T3	I0/I3899/net049	net946	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3899/T4	vss	I0/I3899/net13	I0/I3899/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3899/T5	I0/I3899/net13	I0/I3899/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3899/T2	BL31	net946	I0/I3899/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3867/T3	I0/I3867/net049	net946	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3867/T4	vss	I0/I3867/net13	I0/I3867/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3889/T3	I0/I3889/net049	net945	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3889/T4	vss	I0/I3889/net13	I0/I3889/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3889/T5	I0/I3889/net13	I0/I3889/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3889/T2	BL31	net945	I0/I3889/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3857/T3	I0/I3857/net049	net945	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3857/T4	vss	I0/I3857/net13	I0/I3857/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3915/T3	I0/I3915/net049	net944	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3915/T4	vss	I0/I3915/net13	I0/I3915/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3915/T5	I0/I3915/net13	I0/I3915/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3915/T2	BL31	net944	I0/I3915/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3883/T3	I0/I3883/net049	net944	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3883/T4	vss	I0/I3883/net13	I0/I3883/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3909/T3	I0/I3909/net049	net943	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3909/T4	vss	I0/I3909/net13	I0/I3909/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3909/T5	I0/I3909/net13	I0/I3909/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3909/T2	BL31	net943	I0/I3909/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3877/T3	I0/I3877/net049	net943	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3877/T4	vss	I0/I3877/net13	I0/I3877/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3895/T3	I0/I3895/net049	net942	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3895/T4	vss	I0/I3895/net13	I0/I3895/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3895/T5	I0/I3895/net13	I0/I3895/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3895/T2	BL31	net942	I0/I3895/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3863/T3	I0/I3863/net049	net942	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3863/T4	vss	I0/I3863/net13	I0/I3863/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3888/T3	I0/I3888/net049	net941	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3888/T4	vss	I0/I3888/net13	I0/I3888/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3888/T5	I0/I3888/net13	I0/I3888/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3888/T2	BL31	net941	I0/I3888/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3856/T3	I0/I3856/net049	net941	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3856/T4	vss	I0/I3856/net13	I0/I3856/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3911/T3	I0/I3911/net049	net940	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3911/T4	vss	I0/I3911/net13	I0/I3911/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3911/T5	I0/I3911/net13	I0/I3911/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3911/T2	BL31	net940	I0/I3911/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3879/T3	I0/I3879/net049	net940	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3879/T4	vss	I0/I3879/net13	I0/I3879/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3908/T3	I0/I3908/net049	net939	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3908/T4	vss	I0/I3908/net13	I0/I3908/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3908/T5	I0/I3908/net13	I0/I3908/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3908/T2	BL31	net939	I0/I3908/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3876/T3	I0/I3876/net049	net939	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3876/T4	vss	I0/I3876/net13	I0/I3876/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3886/T3	I0/I3886/net049	net938	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3886/T4	vss	I0/I3886/net13	I0/I3886/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3886/T5	I0/I3886/net13	I0/I3886/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3886/T2	BL31	net938	I0/I3886/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3854/T3	I0/I3854/net049	net938	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3854/T4	vss	I0/I3854/net13	I0/I3854/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3675/T2	BL24	net946	I0/I3675/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3665/T2	BL24	net945	I0/I3665/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3691/T2	BL24	net944	I0/I3691/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3685/T2	BL24	net943	I0/I3685/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3671/T2	BL24	net942	I0/I3671/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3664/T2	BL24	net941	I0/I3664/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3687/T2	BL24	net940	I0/I3687/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3684/T2	BL24	net939	I0/I3684/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3662/T2	BL24	net938	I0/I3662/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3675/T3	I0/I3675/net049	net946	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3665/T3	I0/I3665/net049	net945	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3675/T4	vss	I0/I3675/net13	I0/I3675/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3665/T4	vss	I0/I3665/net13	I0/I3665/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3675/T5	I0/I3675/net13	I0/I3675/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3665/T5	I0/I3665/net13	I0/I3665/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3691/T3	I0/I3691/net049	net944	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3685/T3	I0/I3685/net049	net943	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3691/T4	vss	I0/I3691/net13	I0/I3691/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3685/T4	vss	I0/I3685/net13	I0/I3685/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3691/T5	I0/I3691/net13	I0/I3691/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3685/T5	I0/I3685/net13	I0/I3685/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3671/T3	I0/I3671/net049	net942	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3671/T4	vss	I0/I3671/net13	I0/I3671/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3671/T5	I0/I3671/net13	I0/I3671/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3664/T3	I0/I3664/net049	net941	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3687/T3	I0/I3687/net049	net940	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3664/T4	vss	I0/I3664/net13	I0/I3664/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3687/T4	vss	I0/I3687/net13	I0/I3687/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3664/T5	I0/I3664/net13	I0/I3664/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3687/T5	I0/I3687/net13	I0/I3687/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3684/T3	I0/I3684/net049	net939	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3662/T3	I0/I3662/net049	net938	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3684/T4	vss	I0/I3684/net13	I0/I3684/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3662/T4	vss	I0/I3662/net13	I0/I3662/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3684/T5	I0/I3684/net13	I0/I3684/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3662/T5	I0/I3662/net13	I0/I3662/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3707/T2	BL25	net946	I0/I3707/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3697/T2	BL25	net945	I0/I3697/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3723/T2	BL25	net944	I0/I3723/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3717/T2	BL25	net943	I0/I3717/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3703/T2	BL25	net942	I0/I3703/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3696/T2	BL25	net941	I0/I3696/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3719/T2	BL25	net940	I0/I3719/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3716/T2	BL25	net939	I0/I3716/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3694/T2	BL25	net938	I0/I3694/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3707/T5	I0/I3707/net13	I0/I3707/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3697/T5	I0/I3697/net13	I0/I3697/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3723/T5	I0/I3723/net13	I0/I3723/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3717/T5	I0/I3717/net13	I0/I3717/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3703/T5	I0/I3703/net13	I0/I3703/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3696/T5	I0/I3696/net13	I0/I3696/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3719/T5	I0/I3719/net13	I0/I3719/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3716/T5	I0/I3716/net13	I0/I3716/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3694/T5	I0/I3694/net13	I0/I3694/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3707/T4	vss	I0/I3707/net13	I0/I3707/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3697/T4	vss	I0/I3697/net13	I0/I3697/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3723/T4	vss	I0/I3723/net13	I0/I3723/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3717/T4	vss	I0/I3717/net13	I0/I3717/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3703/T4	vss	I0/I3703/net13	I0/I3703/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3696/T4	vss	I0/I3696/net13	I0/I3696/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3719/T4	vss	I0/I3719/net13	I0/I3719/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3716/T4	vss	I0/I3716/net13	I0/I3716/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3694/T4	vss	I0/I3694/net13	I0/I3694/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3707/T3	I0/I3707/net049	net946	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3697/T3	I0/I3697/net049	net945	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3723/T3	I0/I3723/net049	net944	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3717/T3	I0/I3717/net049	net943	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3703/T3	I0/I3703/net049	net942	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3696/T3	I0/I3696/net049	net941	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3719/T3	I0/I3719/net049	net940	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3716/T3	I0/I3716/net049	net939	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3694/T3	I0/I3694/net049	net938	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3887/T3	I0/I3887/net049	net937	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3887/T4	vss	I0/I3887/net13	I0/I3887/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3887/T5	I0/I3887/net13	I0/I3887/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3887/T2	BL31	net937	I0/I3887/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3855/T3	I0/I3855/net049	net937	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3855/T4	vss	I0/I3855/net13	I0/I3855/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3663/T2	BL24	net937	I0/I3663/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3695/T3	I0/I3695/net049	net937	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3695/T4	vss	I0/I3695/net13	I0/I3695/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3695/T5	I0/I3695/net13	I0/I3695/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3695/T2	BL25	net937	I0/I3695/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3663/T3	I0/I3663/net049	net937	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3663/T4	vss	I0/I3663/net13	I0/I3663/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3663/T5	I0/I3663/net13	I0/I3663/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3894/T3	I0/I3894/net049	net936	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3894/T4	vss	I0/I3894/net13	I0/I3894/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3894/T5	I0/I3894/net13	I0/I3894/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3894/T2	BL31	net936	I0/I3894/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3862/T3	I0/I3862/net049	net936	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3862/T4	vss	I0/I3862/net13	I0/I3862/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3670/T2	BL24	net936	I0/I3670/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3702/T3	I0/I3702/net049	net936	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3702/T4	vss	I0/I3702/net13	I0/I3702/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3702/T5	I0/I3702/net13	I0/I3702/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3702/T2	BL25	net936	I0/I3702/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3670/T3	I0/I3670/net049	net936	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3670/T4	vss	I0/I3670/net13	I0/I3670/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3670/T5	I0/I3670/net13	I0/I3670/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3896/T3	I0/I3896/net049	net935	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3896/T4	vss	I0/I3896/net13	I0/I3896/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3896/T5	I0/I3896/net13	I0/I3896/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3896/T2	BL31	net935	I0/I3896/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3864/T3	I0/I3864/net049	net935	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3864/T4	vss	I0/I3864/net13	I0/I3864/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3672/T2	BL24	net935	I0/I3672/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3704/T3	I0/I3704/net049	net935	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3704/T4	vss	I0/I3704/net13	I0/I3704/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3704/T5	I0/I3704/net13	I0/I3704/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3704/T2	BL25	net935	I0/I3704/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3672/T3	I0/I3672/net049	net935	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3672/T4	vss	I0/I3672/net13	I0/I3672/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3672/T5	I0/I3672/net13	I0/I3672/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3902/T3	I0/I3902/net049	net934	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3902/T4	vss	I0/I3902/net13	I0/I3902/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3902/T5	I0/I3902/net13	I0/I3902/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3902/T2	BL31	net934	I0/I3902/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3870/T3	I0/I3870/net049	net934	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3870/T4	vss	I0/I3870/net13	I0/I3870/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3678/T2	BL24	net934	I0/I3678/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3710/T3	I0/I3710/net049	net934	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3710/T4	vss	I0/I3710/net13	I0/I3710/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3710/T5	I0/I3710/net13	I0/I3710/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3710/T2	BL25	net934	I0/I3710/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3678/T3	I0/I3678/net049	net934	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3678/T4	vss	I0/I3678/net13	I0/I3678/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3678/T5	I0/I3678/net13	I0/I3678/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3904/T3	I0/I3904/net049	net933	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3904/T4	vss	I0/I3904/net13	I0/I3904/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3904/T5	I0/I3904/net13	I0/I3904/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3904/T2	BL31	net933	I0/I3904/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3872/T3	I0/I3872/net049	net933	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3872/T4	vss	I0/I3872/net13	I0/I3872/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3680/T2	BL24	net933	I0/I3680/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3712/T3	I0/I3712/net049	net933	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3712/T4	vss	I0/I3712/net13	I0/I3712/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3712/T5	I0/I3712/net13	I0/I3712/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3712/T2	BL25	net933	I0/I3712/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3680/T3	I0/I3680/net049	net933	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3680/T4	vss	I0/I3680/net13	I0/I3680/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3680/T5	I0/I3680/net13	I0/I3680/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3893/T3	I0/I3893/net049	net932	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3893/T4	vss	I0/I3893/net13	I0/I3893/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3893/T5	I0/I3893/net13	I0/I3893/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3893/T2	BL31	net932	I0/I3893/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3861/T3	I0/I3861/net049	net932	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3861/T4	vss	I0/I3861/net13	I0/I3861/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3669/T2	BL24	net932	I0/I3669/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3701/T3	I0/I3701/net049	net932	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3701/T4	vss	I0/I3701/net13	I0/I3701/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3701/T5	I0/I3701/net13	I0/I3701/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3701/T2	BL25	net932	I0/I3701/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3669/T3	I0/I3669/net049	net932	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3669/T4	vss	I0/I3669/net13	I0/I3669/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3669/T5	I0/I3669/net13	I0/I3669/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3907/T3	I0/I3907/net049	net931	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3907/T4	vss	I0/I3907/net13	I0/I3907/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3907/T5	I0/I3907/net13	I0/I3907/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3907/T2	BL31	net931	I0/I3907/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3875/T3	I0/I3875/net049	net931	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3875/T4	vss	I0/I3875/net13	I0/I3875/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3683/T2	BL24	net931	I0/I3683/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3715/T3	I0/I3715/net049	net931	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3715/T4	vss	I0/I3715/net13	I0/I3715/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3715/T5	I0/I3715/net13	I0/I3715/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3715/T2	BL25	net931	I0/I3715/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3683/T3	I0/I3683/net049	net931	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3683/T4	vss	I0/I3683/net13	I0/I3683/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3683/T5	I0/I3683/net13	I0/I3683/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3901/T3	I0/I3901/net049	net930	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3901/T4	vss	I0/I3901/net13	I0/I3901/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3901/T5	I0/I3901/net13	I0/I3901/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3901/T2	BL31	net930	I0/I3901/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3869/T3	I0/I3869/net049	net930	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3869/T4	vss	I0/I3869/net13	I0/I3869/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3677/T2	BL24	net930	I0/I3677/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3709/T3	I0/I3709/net049	net930	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3709/T4	vss	I0/I3709/net13	I0/I3709/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3709/T5	I0/I3709/net13	I0/I3709/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3709/T2	BL25	net930	I0/I3709/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3677/T3	I0/I3677/net049	net930	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3677/T4	vss	I0/I3677/net13	I0/I3677/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3677/T5	I0/I3677/net13	I0/I3677/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3905/T3	I0/I3905/net049	net929	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3905/T4	vss	I0/I3905/net13	I0/I3905/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3905/T5	I0/I3905/net13	I0/I3905/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3905/T2	BL31	net929	I0/I3905/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3873/T3	I0/I3873/net049	net929	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3873/T4	vss	I0/I3873/net13	I0/I3873/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3681/T2	BL24	net929	I0/I3681/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3713/T3	I0/I3713/net049	net929	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3713/T4	vss	I0/I3713/net13	I0/I3713/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3713/T5	I0/I3713/net13	I0/I3713/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3713/T2	BL25	net929	I0/I3713/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3681/T3	I0/I3681/net049	net929	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3681/T4	vss	I0/I3681/net13	I0/I3681/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3681/T5	I0/I3681/net13	I0/I3681/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3917/T3	I0/I3917/net049	net928	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3917/T4	vss	I0/I3917/net13	I0/I3917/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3917/T5	I0/I3917/net13	I0/I3917/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3917/T2	BL31	net928	I0/I3917/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3885/T3	I0/I3885/net049	net928	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3885/T4	vss	I0/I3885/net13	I0/I3885/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3693/T2	BL24	net928	I0/I3693/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3725/T3	I0/I3725/net049	net928	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3725/T4	vss	I0/I3725/net13	I0/I3725/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3725/T5	I0/I3725/net13	I0/I3725/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3725/T2	BL25	net928	I0/I3725/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3693/T3	I0/I3693/net049	net928	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3693/T4	vss	I0/I3693/net13	I0/I3693/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3693/T5	I0/I3693/net13	I0/I3693/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3903/T3	I0/I3903/net049	net927	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3903/T4	vss	I0/I3903/net13	I0/I3903/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3903/T5	I0/I3903/net13	I0/I3903/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3903/T2	BL31	net927	I0/I3903/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3871/T3	I0/I3871/net049	net927	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3871/T4	vss	I0/I3871/net13	I0/I3871/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3679/T2	BL24	net927	I0/I3679/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3711/T3	I0/I3711/net049	net927	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3711/T4	vss	I0/I3711/net13	I0/I3711/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3711/T5	I0/I3711/net13	I0/I3711/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3711/T2	BL25	net927	I0/I3711/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3679/T3	I0/I3679/net049	net927	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3679/T4	vss	I0/I3679/net13	I0/I3679/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3679/T5	I0/I3679/net13	I0/I3679/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3914/T3	I0/I3914/net049	net926	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3914/T4	vss	I0/I3914/net13	I0/I3914/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3914/T5	I0/I3914/net13	I0/I3914/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3914/T2	BL31	net926	I0/I3914/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3882/T3	I0/I3882/net049	net926	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3882/T4	vss	I0/I3882/net13	I0/I3882/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3690/T2	BL24	net926	I0/I3690/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3722/T3	I0/I3722/net049	net926	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3722/T4	vss	I0/I3722/net13	I0/I3722/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3722/T5	I0/I3722/net13	I0/I3722/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3722/T2	BL25	net926	I0/I3722/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3690/T3	I0/I3690/net049	net926	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3690/T4	vss	I0/I3690/net13	I0/I3690/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3690/T5	I0/I3690/net13	I0/I3690/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3913/T3	I0/I3913/net049	net925	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3913/T4	vss	I0/I3913/net13	I0/I3913/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3913/T5	I0/I3913/net13	I0/I3913/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3913/T2	BL31	net925	I0/I3913/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3881/T3	I0/I3881/net049	net925	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3881/T4	vss	I0/I3881/net13	I0/I3881/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3689/T2	BL24	net925	I0/I3689/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3721/T3	I0/I3721/net049	net925	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3721/T4	vss	I0/I3721/net13	I0/I3721/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3721/T5	I0/I3721/net13	I0/I3721/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3721/T2	BL25	net925	I0/I3721/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3689/T3	I0/I3689/net049	net925	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3689/T4	vss	I0/I3689/net13	I0/I3689/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3689/T5	I0/I3689/net13	I0/I3689/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3890/T3	I0/I3890/net049	net924	BL31bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3890/T4	vss	I0/I3890/net13	I0/I3890/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3890/T5	I0/I3890/net13	I0/I3890/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3890/T2	BL31	net924	I0/I3890/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3858/T3	I0/I3858/net049	net924	BL30bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3858/T4	vss	I0/I3858/net13	I0/I3858/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3666/T2	BL24	net924	I0/I3666/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3698/T3	I0/I3698/net049	net924	BL25bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3698/T4	vss	I0/I3698/net13	I0/I3698/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3698/T5	I0/I3698/net13	I0/I3698/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3698/T2	BL25	net924	I0/I3698/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3666/T3	I0/I3666/net049	net924	BL24bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3666/T4	vss	I0/I3666/net13	I0/I3666/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3666/T5	I0/I3666/net13	I0/I3666/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI88/T1	p7bar	y2	BL25bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI89/T1	BL25	y2	p7	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI90/T1	p7bar	y1	BL24bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI91/T1	BL24	y1	p7	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI92/T1	p8bar	y4	BL31bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI93/T1	BL31	y4	p8	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI94/T1	p8bar	y3	BL30bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T8	vss	I6/net20	I6/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T7	data5	I6/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T11	I28/net23	data5	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T16	I28/net15	net680	p6	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T17	vss	I28/net23	I28/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T19	I28/net7	p6	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T18	p6bar	net680	I28/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T2	I7/net23	p7	I7/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T3	I7/net20	p7bar	I7/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T4	vss	vdd	I7/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T8	vss	I7/net20	I7/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T7	data6	I7/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3740/T2	BL26	net955	I0/I3740/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3732/T2	BL26	net954	I0/I3732/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3731/T2	BL26	net953	I0/I3731/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3756/T2	BL26	net952	I0/I3756/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3737/T2	BL26	net951	I0/I3737/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3752/T2	BL26	net950	I0/I3752/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3750/T2	BL26	net949	I0/I3750/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3746/T2	BL26	net948	I0/I3746/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3738/T2	BL26	net947	I0/I3738/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3739/T2	BL26	net946	I0/I3739/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3729/T2	BL26	net945	I0/I3729/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3755/T2	BL26	net944	I0/I3755/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3749/T2	BL26	net943	I0/I3749/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3735/T2	BL26	net942	I0/I3735/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3728/T2	BL26	net941	I0/I3728/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3751/T2	BL26	net940	I0/I3751/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3748/T2	BL26	net939	I0/I3748/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3726/T2	BL26	net938	I0/I3726/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3727/T2	BL26	net937	I0/I3727/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3734/T2	BL26	net936	I0/I3734/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3736/T2	BL26	net935	I0/I3736/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3742/T2	BL26	net934	I0/I3742/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3744/T2	BL26	net933	I0/I3744/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3733/T2	BL26	net932	I0/I3733/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3747/T2	BL26	net931	I0/I3747/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3741/T2	BL26	net930	I0/I3741/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3745/T2	BL26	net929	I0/I3745/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3757/T2	BL26	net928	I0/I3757/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3743/T2	BL26	net927	I0/I3743/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3754/T2	BL26	net926	I0/I3754/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3753/T2	BL26	net925	I0/I3753/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3730/T2	BL26	net924	I0/I3730/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI87/T1	BL26	y3	p7	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T4	vss	vdd	I6/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3740/T3	I0/I3740/net049	net955	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3732/T3	I0/I3732/net049	net954	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3740/T4	vss	I0/I3740/net13	I0/I3740/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3732/T4	vss	I0/I3732/net13	I0/I3732/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3740/T5	I0/I3740/net13	I0/I3740/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3732/T5	I0/I3732/net13	I0/I3732/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3731/T3	I0/I3731/net049	net953	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3756/T3	I0/I3756/net049	net952	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3731/T4	vss	I0/I3731/net13	I0/I3731/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3756/T4	vss	I0/I3756/net13	I0/I3756/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3731/T5	I0/I3731/net13	I0/I3731/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3756/T5	I0/I3756/net13	I0/I3756/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3737/T3	I0/I3737/net049	net951	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3737/T4	vss	I0/I3737/net13	I0/I3737/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3737/T5	I0/I3737/net13	I0/I3737/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3752/T3	I0/I3752/net049	net950	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3750/T3	I0/I3750/net049	net949	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3752/T4	vss	I0/I3752/net13	I0/I3752/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3750/T4	vss	I0/I3750/net13	I0/I3750/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3752/T5	I0/I3752/net13	I0/I3752/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3750/T5	I0/I3750/net13	I0/I3750/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3746/T3	I0/I3746/net049	net948	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3738/T3	I0/I3738/net049	net947	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3746/T4	vss	I0/I3746/net13	I0/I3746/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3738/T4	vss	I0/I3738/net13	I0/I3738/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3746/T5	I0/I3746/net13	I0/I3746/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3738/T5	I0/I3738/net13	I0/I3738/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3772/T2	BL27	net955	I0/I3772/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3764/T2	BL27	net954	I0/I3764/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3763/T2	BL27	net953	I0/I3763/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3788/T2	BL27	net952	I0/I3788/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3769/T2	BL27	net951	I0/I3769/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3784/T2	BL27	net950	I0/I3784/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3782/T2	BL27	net949	I0/I3782/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3778/T2	BL27	net948	I0/I3778/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3770/T2	BL27	net947	I0/I3770/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3772/T5	I0/I3772/net13	I0/I3772/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3764/T5	I0/I3764/net13	I0/I3764/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3763/T5	I0/I3763/net13	I0/I3763/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3788/T5	I0/I3788/net13	I0/I3788/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3769/T5	I0/I3769/net13	I0/I3769/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3784/T5	I0/I3784/net13	I0/I3784/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3782/T5	I0/I3782/net13	I0/I3782/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3778/T5	I0/I3778/net13	I0/I3778/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3770/T5	I0/I3770/net13	I0/I3770/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3772/T4	vss	I0/I3772/net13	I0/I3772/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3764/T4	vss	I0/I3764/net13	I0/I3764/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3763/T4	vss	I0/I3763/net13	I0/I3763/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3788/T4	vss	I0/I3788/net13	I0/I3788/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3769/T4	vss	I0/I3769/net13	I0/I3769/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3784/T4	vss	I0/I3784/net13	I0/I3784/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3782/T4	vss	I0/I3782/net13	I0/I3782/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3778/T4	vss	I0/I3778/net13	I0/I3778/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3770/T4	vss	I0/I3770/net13	I0/I3770/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3772/T3	I0/I3772/net049	net955	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3764/T3	I0/I3764/net049	net954	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3763/T3	I0/I3763/net049	net953	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3788/T3	I0/I3788/net049	net952	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3769/T3	I0/I3769/net049	net951	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3784/T3	I0/I3784/net049	net950	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3782/T3	I0/I3782/net049	net949	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3778/T3	I0/I3778/net049	net948	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3770/T3	I0/I3770/net049	net947	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3548/T2	BL20	net955	I0/I3548/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3540/T2	BL20	net954	I0/I3540/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3539/T2	BL20	net953	I0/I3539/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3564/T2	BL20	net952	I0/I3564/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3545/T2	BL20	net951	I0/I3545/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3560/T2	BL20	net950	I0/I3560/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3558/T2	BL20	net949	I0/I3558/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3554/T2	BL20	net948	I0/I3554/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3546/T2	BL20	net947	I0/I3546/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3548/T5	I0/I3548/net13	I0/I3548/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3540/T5	I0/I3540/net13	I0/I3540/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3539/T5	I0/I3539/net13	I0/I3539/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3564/T5	I0/I3564/net13	I0/I3564/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3545/T5	I0/I3545/net13	I0/I3545/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3560/T5	I0/I3560/net13	I0/I3560/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3558/T5	I0/I3558/net13	I0/I3558/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3554/T5	I0/I3554/net13	I0/I3554/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3546/T5	I0/I3546/net13	I0/I3546/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3548/T4	vss	I0/I3548/net13	I0/I3548/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3540/T4	vss	I0/I3540/net13	I0/I3540/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3539/T4	vss	I0/I3539/net13	I0/I3539/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3564/T4	vss	I0/I3564/net13	I0/I3564/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3545/T4	vss	I0/I3545/net13	I0/I3545/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3560/T4	vss	I0/I3560/net13	I0/I3560/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3558/T4	vss	I0/I3558/net13	I0/I3558/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3554/T4	vss	I0/I3554/net13	I0/I3554/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3546/T4	vss	I0/I3546/net13	I0/I3546/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3548/T3	I0/I3548/net049	net955	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3540/T3	I0/I3540/net049	net954	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3539/T3	I0/I3539/net049	net953	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3564/T3	I0/I3564/net049	net952	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3545/T3	I0/I3545/net049	net951	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3560/T3	I0/I3560/net049	net950	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3558/T3	I0/I3558/net049	net949	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3554/T3	I0/I3554/net049	net948	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3546/T3	I0/I3546/net049	net947	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3580/T4	vss	I0/I3580/net13	I0/I3580/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3572/T4	vss	I0/I3572/net13	I0/I3572/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3580/T5	I0/I3580/net13	I0/I3580/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3572/T5	I0/I3572/net13	I0/I3572/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3580/T2	BL21	net955	I0/I3580/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3572/T2	BL21	net954	I0/I3572/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3571/T4	vss	I0/I3571/net13	I0/I3571/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3596/T4	vss	I0/I3596/net13	I0/I3596/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3571/T5	I0/I3571/net13	I0/I3571/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3596/T5	I0/I3596/net13	I0/I3596/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3571/T2	BL21	net953	I0/I3571/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3596/T2	BL21	net952	I0/I3596/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3577/T4	vss	I0/I3577/net13	I0/I3577/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3577/T5	I0/I3577/net13	I0/I3577/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3577/T2	BL21	net951	I0/I3577/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3592/T4	vss	I0/I3592/net13	I0/I3592/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3590/T4	vss	I0/I3590/net13	I0/I3590/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3592/T5	I0/I3592/net13	I0/I3592/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3590/T5	I0/I3590/net13	I0/I3590/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3592/T2	BL21	net950	I0/I3592/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3590/T2	BL21	net949	I0/I3590/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3586/T4	vss	I0/I3586/net13	I0/I3586/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3578/T4	vss	I0/I3578/net13	I0/I3578/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3586/T5	I0/I3586/net13	I0/I3586/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3578/T5	I0/I3578/net13	I0/I3578/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3586/T2	BL21	net948	I0/I3586/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3578/T2	BL21	net947	I0/I3578/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3580/T3	I0/I3580/net049	net955	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3572/T3	I0/I3572/net049	net954	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3571/T3	I0/I3571/net049	net953	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3596/T3	I0/I3596/net049	net952	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3577/T3	I0/I3577/net049	net951	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3592/T3	I0/I3592/net049	net950	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3590/T3	I0/I3590/net049	net949	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3586/T3	I0/I3586/net049	net948	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3578/T3	I0/I3578/net049	net947	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3612/T2	BL22	net955	I0/I3612/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3604/T2	BL22	net954	I0/I3604/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3603/T2	BL22	net953	I0/I3603/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3628/T2	BL22	net952	I0/I3628/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3609/T2	BL22	net951	I0/I3609/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3624/T2	BL22	net950	I0/I3624/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3622/T2	BL22	net949	I0/I3622/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3618/T2	BL22	net948	I0/I3618/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3610/T2	BL22	net947	I0/I3610/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3612/T5	I0/I3612/net13	I0/I3612/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3604/T5	I0/I3604/net13	I0/I3604/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3603/T5	I0/I3603/net13	I0/I3603/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3628/T5	I0/I3628/net13	I0/I3628/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3609/T5	I0/I3609/net13	I0/I3609/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3624/T5	I0/I3624/net13	I0/I3624/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3622/T5	I0/I3622/net13	I0/I3622/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3618/T5	I0/I3618/net13	I0/I3618/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3610/T5	I0/I3610/net13	I0/I3610/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3612/T4	vss	I0/I3612/net13	I0/I3612/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3604/T4	vss	I0/I3604/net13	I0/I3604/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3603/T4	vss	I0/I3603/net13	I0/I3603/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3628/T4	vss	I0/I3628/net13	I0/I3628/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3609/T4	vss	I0/I3609/net13	I0/I3609/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3624/T4	vss	I0/I3624/net13	I0/I3624/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3622/T4	vss	I0/I3622/net13	I0/I3622/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3618/T4	vss	I0/I3618/net13	I0/I3618/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3610/T4	vss	I0/I3610/net13	I0/I3610/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3612/T3	I0/I3612/net049	net955	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3604/T3	I0/I3604/net049	net954	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3603/T3	I0/I3603/net049	net953	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3628/T3	I0/I3628/net049	net952	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3609/T3	I0/I3609/net049	net951	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3624/T3	I0/I3624/net049	net950	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3622/T3	I0/I3622/net049	net949	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3618/T3	I0/I3618/net049	net948	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3610/T3	I0/I3610/net049	net947	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3644/T4	vss	I0/I3644/net13	I0/I3644/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3636/T4	vss	I0/I3636/net13	I0/I3636/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3644/T5	I0/I3644/net13	I0/I3644/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3636/T5	I0/I3636/net13	I0/I3636/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3644/T2	BL23	net955	I0/I3644/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3636/T2	BL23	net954	I0/I3636/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3635/T4	vss	I0/I3635/net13	I0/I3635/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3660/T4	vss	I0/I3660/net13	I0/I3660/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3635/T5	I0/I3635/net13	I0/I3635/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3660/T5	I0/I3660/net13	I0/I3660/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3635/T2	BL23	net953	I0/I3635/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3660/T2	BL23	net952	I0/I3660/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3641/T4	vss	I0/I3641/net13	I0/I3641/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3641/T5	I0/I3641/net13	I0/I3641/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3641/T2	BL23	net951	I0/I3641/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3656/T4	vss	I0/I3656/net13	I0/I3656/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3654/T4	vss	I0/I3654/net13	I0/I3654/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3656/T5	I0/I3656/net13	I0/I3656/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3654/T5	I0/I3654/net13	I0/I3654/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3656/T2	BL23	net950	I0/I3656/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3654/T2	BL23	net949	I0/I3654/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3650/T4	vss	I0/I3650/net13	I0/I3650/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3642/T4	vss	I0/I3642/net13	I0/I3642/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3650/T5	I0/I3650/net13	I0/I3650/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3642/T5	I0/I3642/net13	I0/I3642/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3650/T2	BL23	net948	I0/I3650/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3642/T2	BL23	net947	I0/I3642/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3644/T3	I0/I3644/net049	net955	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3636/T3	I0/I3636/net049	net954	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3635/T3	I0/I3635/net049	net953	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3660/T3	I0/I3660/net049	net952	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3641/T3	I0/I3641/net049	net951	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3656/T3	I0/I3656/net049	net950	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3654/T3	I0/I3654/net049	net949	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3650/T3	I0/I3650/net049	net948	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3642/T3	I0/I3642/net049	net947	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3420/T2	BL16	net955	I0/I3420/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3412/T2	BL16	net954	I0/I3412/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3411/T2	BL16	net953	I0/I3411/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3436/T2	BL16	net952	I0/I3436/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3417/T2	BL16	net951	I0/I3417/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3432/T2	BL16	net950	I0/I3432/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3430/T2	BL16	net949	I0/I3430/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3426/T2	BL16	net948	I0/I3426/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3418/T2	BL16	net947	I0/I3418/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3420/T5	I0/I3420/net13	I0/I3420/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3412/T5	I0/I3412/net13	I0/I3412/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3411/T5	I0/I3411/net13	I0/I3411/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3436/T5	I0/I3436/net13	I0/I3436/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3417/T5	I0/I3417/net13	I0/I3417/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3432/T5	I0/I3432/net13	I0/I3432/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3430/T5	I0/I3430/net13	I0/I3430/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3426/T5	I0/I3426/net13	I0/I3426/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3418/T5	I0/I3418/net13	I0/I3418/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3420/T4	vss	I0/I3420/net13	I0/I3420/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3412/T4	vss	I0/I3412/net13	I0/I3412/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3411/T4	vss	I0/I3411/net13	I0/I3411/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3436/T4	vss	I0/I3436/net13	I0/I3436/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3417/T4	vss	I0/I3417/net13	I0/I3417/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3432/T4	vss	I0/I3432/net13	I0/I3432/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3430/T4	vss	I0/I3430/net13	I0/I3430/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3426/T4	vss	I0/I3426/net13	I0/I3426/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3418/T4	vss	I0/I3418/net13	I0/I3418/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3420/T3	I0/I3420/net049	net955	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3412/T3	I0/I3412/net049	net954	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3411/T3	I0/I3411/net049	net953	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3436/T3	I0/I3436/net049	net952	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3417/T3	I0/I3417/net049	net951	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3432/T3	I0/I3432/net049	net950	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3430/T3	I0/I3430/net049	net949	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3426/T3	I0/I3426/net049	net948	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3418/T3	I0/I3418/net049	net947	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3452/T2	BL17	net955	I0/I3452/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3444/T2	BL17	net954	I0/I3444/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3443/T2	BL17	net953	I0/I3443/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3468/T2	BL17	net952	I0/I3468/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3449/T2	BL17	net951	I0/I3449/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3464/T2	BL17	net950	I0/I3464/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3462/T2	BL17	net949	I0/I3462/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3458/T2	BL17	net948	I0/I3458/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3450/T2	BL17	net947	I0/I3450/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3739/T3	I0/I3739/net049	net946	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3729/T3	I0/I3729/net049	net945	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3739/T4	vss	I0/I3739/net13	I0/I3739/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3729/T4	vss	I0/I3729/net13	I0/I3729/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3739/T5	I0/I3739/net13	I0/I3739/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3729/T5	I0/I3729/net13	I0/I3729/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3755/T3	I0/I3755/net049	net944	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3749/T3	I0/I3749/net049	net943	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3755/T4	vss	I0/I3755/net13	I0/I3755/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3749/T4	vss	I0/I3749/net13	I0/I3749/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3755/T5	I0/I3755/net13	I0/I3755/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3749/T5	I0/I3749/net13	I0/I3749/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3735/T3	I0/I3735/net049	net942	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3735/T4	vss	I0/I3735/net13	I0/I3735/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3735/T5	I0/I3735/net13	I0/I3735/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3728/T3	I0/I3728/net049	net941	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3751/T3	I0/I3751/net049	net940	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3728/T4	vss	I0/I3728/net13	I0/I3728/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3751/T4	vss	I0/I3751/net13	I0/I3751/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3728/T5	I0/I3728/net13	I0/I3728/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3751/T5	I0/I3751/net13	I0/I3751/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3748/T3	I0/I3748/net049	net939	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3726/T3	I0/I3726/net049	net938	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3748/T4	vss	I0/I3748/net13	I0/I3748/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3726/T4	vss	I0/I3726/net13	I0/I3726/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3748/T5	I0/I3748/net13	I0/I3748/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3726/T5	I0/I3726/net13	I0/I3726/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3771/T2	BL27	net946	I0/I3771/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3761/T2	BL27	net945	I0/I3761/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3787/T2	BL27	net944	I0/I3787/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3781/T2	BL27	net943	I0/I3781/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3767/T2	BL27	net942	I0/I3767/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3760/T2	BL27	net941	I0/I3760/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3783/T2	BL27	net940	I0/I3783/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3780/T2	BL27	net939	I0/I3780/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3758/T2	BL27	net938	I0/I3758/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3771/T5	I0/I3771/net13	I0/I3771/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3761/T5	I0/I3761/net13	I0/I3761/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3787/T5	I0/I3787/net13	I0/I3787/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3781/T5	I0/I3781/net13	I0/I3781/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3767/T5	I0/I3767/net13	I0/I3767/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3760/T5	I0/I3760/net13	I0/I3760/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3783/T5	I0/I3783/net13	I0/I3783/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3780/T5	I0/I3780/net13	I0/I3780/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3758/T5	I0/I3758/net13	I0/I3758/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3771/T4	vss	I0/I3771/net13	I0/I3771/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3761/T4	vss	I0/I3761/net13	I0/I3761/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3787/T4	vss	I0/I3787/net13	I0/I3787/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3781/T4	vss	I0/I3781/net13	I0/I3781/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3767/T4	vss	I0/I3767/net13	I0/I3767/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3760/T4	vss	I0/I3760/net13	I0/I3760/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3783/T4	vss	I0/I3783/net13	I0/I3783/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3780/T4	vss	I0/I3780/net13	I0/I3780/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3758/T4	vss	I0/I3758/net13	I0/I3758/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3771/T3	I0/I3771/net049	net946	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3761/T3	I0/I3761/net049	net945	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3787/T3	I0/I3787/net049	net944	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3781/T3	I0/I3781/net049	net943	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3767/T3	I0/I3767/net049	net942	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3760/T3	I0/I3760/net049	net941	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3783/T3	I0/I3783/net049	net940	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3780/T3	I0/I3780/net049	net939	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3758/T3	I0/I3758/net049	net938	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3547/T2	BL20	net946	I0/I3547/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3537/T2	BL20	net945	I0/I3537/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3563/T2	BL20	net944	I0/I3563/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3557/T2	BL20	net943	I0/I3557/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3543/T2	BL20	net942	I0/I3543/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3536/T2	BL20	net941	I0/I3536/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3559/T2	BL20	net940	I0/I3559/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3556/T2	BL20	net939	I0/I3556/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3534/T2	BL20	net938	I0/I3534/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3547/T5	I0/I3547/net13	I0/I3547/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3537/T5	I0/I3537/net13	I0/I3537/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3563/T5	I0/I3563/net13	I0/I3563/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3557/T5	I0/I3557/net13	I0/I3557/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3543/T5	I0/I3543/net13	I0/I3543/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3536/T5	I0/I3536/net13	I0/I3536/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3559/T5	I0/I3559/net13	I0/I3559/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3556/T5	I0/I3556/net13	I0/I3556/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3534/T5	I0/I3534/net13	I0/I3534/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3547/T4	vss	I0/I3547/net13	I0/I3547/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3537/T4	vss	I0/I3537/net13	I0/I3537/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3563/T4	vss	I0/I3563/net13	I0/I3563/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3557/T4	vss	I0/I3557/net13	I0/I3557/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3543/T4	vss	I0/I3543/net13	I0/I3543/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3536/T4	vss	I0/I3536/net13	I0/I3536/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3559/T4	vss	I0/I3559/net13	I0/I3559/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3556/T4	vss	I0/I3556/net13	I0/I3556/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3534/T4	vss	I0/I3534/net13	I0/I3534/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3547/T3	I0/I3547/net049	net946	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3537/T3	I0/I3537/net049	net945	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3563/T3	I0/I3563/net049	net944	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3557/T3	I0/I3557/net049	net943	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3543/T3	I0/I3543/net049	net942	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3536/T3	I0/I3536/net049	net941	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3559/T3	I0/I3559/net049	net940	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3556/T3	I0/I3556/net049	net939	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3534/T3	I0/I3534/net049	net938	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3579/T4	vss	I0/I3579/net13	I0/I3579/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3569/T4	vss	I0/I3569/net13	I0/I3569/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3579/T5	I0/I3579/net13	I0/I3579/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3569/T5	I0/I3569/net13	I0/I3569/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3579/T2	BL21	net946	I0/I3579/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3569/T2	BL21	net945	I0/I3569/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3595/T4	vss	I0/I3595/net13	I0/I3595/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3589/T4	vss	I0/I3589/net13	I0/I3589/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3595/T5	I0/I3595/net13	I0/I3595/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3589/T5	I0/I3589/net13	I0/I3589/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3595/T2	BL21	net944	I0/I3595/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3589/T2	BL21	net943	I0/I3589/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3575/T4	vss	I0/I3575/net13	I0/I3575/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3575/T5	I0/I3575/net13	I0/I3575/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3575/T2	BL21	net942	I0/I3575/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3568/T4	vss	I0/I3568/net13	I0/I3568/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3591/T4	vss	I0/I3591/net13	I0/I3591/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3568/T5	I0/I3568/net13	I0/I3568/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3591/T5	I0/I3591/net13	I0/I3591/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3568/T2	BL21	net941	I0/I3568/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3591/T2	BL21	net940	I0/I3591/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3588/T4	vss	I0/I3588/net13	I0/I3588/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3566/T4	vss	I0/I3566/net13	I0/I3566/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3588/T5	I0/I3588/net13	I0/I3588/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3566/T5	I0/I3566/net13	I0/I3566/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3588/T2	BL21	net939	I0/I3588/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3566/T2	BL21	net938	I0/I3566/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3579/T3	I0/I3579/net049	net946	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3569/T3	I0/I3569/net049	net945	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3595/T3	I0/I3595/net049	net944	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3589/T3	I0/I3589/net049	net943	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3575/T3	I0/I3575/net049	net942	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3568/T3	I0/I3568/net049	net941	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3591/T3	I0/I3591/net049	net940	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3588/T3	I0/I3588/net049	net939	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3566/T3	I0/I3566/net049	net938	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3611/T2	BL22	net946	I0/I3611/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3601/T2	BL22	net945	I0/I3601/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3627/T2	BL22	net944	I0/I3627/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3621/T2	BL22	net943	I0/I3621/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3607/T2	BL22	net942	I0/I3607/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3600/T2	BL22	net941	I0/I3600/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3623/T2	BL22	net940	I0/I3623/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3620/T2	BL22	net939	I0/I3620/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3598/T2	BL22	net938	I0/I3598/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3611/T5	I0/I3611/net13	I0/I3611/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3601/T5	I0/I3601/net13	I0/I3601/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3627/T5	I0/I3627/net13	I0/I3627/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3621/T5	I0/I3621/net13	I0/I3621/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3607/T5	I0/I3607/net13	I0/I3607/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3600/T5	I0/I3600/net13	I0/I3600/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3623/T5	I0/I3623/net13	I0/I3623/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3620/T5	I0/I3620/net13	I0/I3620/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3598/T5	I0/I3598/net13	I0/I3598/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3611/T4	vss	I0/I3611/net13	I0/I3611/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3601/T4	vss	I0/I3601/net13	I0/I3601/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3627/T4	vss	I0/I3627/net13	I0/I3627/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3621/T4	vss	I0/I3621/net13	I0/I3621/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3607/T4	vss	I0/I3607/net13	I0/I3607/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3600/T4	vss	I0/I3600/net13	I0/I3600/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3623/T4	vss	I0/I3623/net13	I0/I3623/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3620/T4	vss	I0/I3620/net13	I0/I3620/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3598/T4	vss	I0/I3598/net13	I0/I3598/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3611/T3	I0/I3611/net049	net946	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3601/T3	I0/I3601/net049	net945	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3627/T3	I0/I3627/net049	net944	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3621/T3	I0/I3621/net049	net943	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3607/T3	I0/I3607/net049	net942	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3600/T3	I0/I3600/net049	net941	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3623/T3	I0/I3623/net049	net940	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3620/T3	I0/I3620/net049	net939	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3598/T3	I0/I3598/net049	net938	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3643/T4	vss	I0/I3643/net13	I0/I3643/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3633/T4	vss	I0/I3633/net13	I0/I3633/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3643/T5	I0/I3643/net13	I0/I3643/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3633/T5	I0/I3633/net13	I0/I3633/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3643/T2	BL23	net946	I0/I3643/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3633/T2	BL23	net945	I0/I3633/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3659/T4	vss	I0/I3659/net13	I0/I3659/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3653/T4	vss	I0/I3653/net13	I0/I3653/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3659/T5	I0/I3659/net13	I0/I3659/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3653/T5	I0/I3653/net13	I0/I3653/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3659/T2	BL23	net944	I0/I3659/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3653/T2	BL23	net943	I0/I3653/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3639/T4	vss	I0/I3639/net13	I0/I3639/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3639/T5	I0/I3639/net13	I0/I3639/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3639/T2	BL23	net942	I0/I3639/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3632/T4	vss	I0/I3632/net13	I0/I3632/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3655/T4	vss	I0/I3655/net13	I0/I3655/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3632/T5	I0/I3632/net13	I0/I3632/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3655/T5	I0/I3655/net13	I0/I3655/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3632/T2	BL23	net941	I0/I3632/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3655/T2	BL23	net940	I0/I3655/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3652/T4	vss	I0/I3652/net13	I0/I3652/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3630/T4	vss	I0/I3630/net13	I0/I3630/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3652/T5	I0/I3652/net13	I0/I3652/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3630/T5	I0/I3630/net13	I0/I3630/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3652/T2	BL23	net939	I0/I3652/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3630/T2	BL23	net938	I0/I3630/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3643/T3	I0/I3643/net049	net946	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3633/T3	I0/I3633/net049	net945	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3659/T3	I0/I3659/net049	net944	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3653/T3	I0/I3653/net049	net943	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3639/T3	I0/I3639/net049	net942	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3632/T3	I0/I3632/net049	net941	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3655/T3	I0/I3655/net049	net940	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3652/T3	I0/I3652/net049	net939	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3630/T3	I0/I3630/net049	net938	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3419/T2	BL16	net946	I0/I3419/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3409/T2	BL16	net945	I0/I3409/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3435/T2	BL16	net944	I0/I3435/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3429/T2	BL16	net943	I0/I3429/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3415/T2	BL16	net942	I0/I3415/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3408/T2	BL16	net941	I0/I3408/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3431/T2	BL16	net940	I0/I3431/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3428/T2	BL16	net939	I0/I3428/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3406/T2	BL16	net938	I0/I3406/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3419/T5	I0/I3419/net13	I0/I3419/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3409/T5	I0/I3409/net13	I0/I3409/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3435/T5	I0/I3435/net13	I0/I3435/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3429/T5	I0/I3429/net13	I0/I3429/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3415/T5	I0/I3415/net13	I0/I3415/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3408/T5	I0/I3408/net13	I0/I3408/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3431/T5	I0/I3431/net13	I0/I3431/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3428/T5	I0/I3428/net13	I0/I3428/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3406/T5	I0/I3406/net13	I0/I3406/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3419/T4	vss	I0/I3419/net13	I0/I3419/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3409/T4	vss	I0/I3409/net13	I0/I3409/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3435/T4	vss	I0/I3435/net13	I0/I3435/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3429/T4	vss	I0/I3429/net13	I0/I3429/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3415/T4	vss	I0/I3415/net13	I0/I3415/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3408/T4	vss	I0/I3408/net13	I0/I3408/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3431/T4	vss	I0/I3431/net13	I0/I3431/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3428/T4	vss	I0/I3428/net13	I0/I3428/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3406/T4	vss	I0/I3406/net13	I0/I3406/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3419/T3	I0/I3419/net049	net946	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3409/T3	I0/I3409/net049	net945	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3435/T3	I0/I3435/net049	net944	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3429/T3	I0/I3429/net049	net943	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3415/T3	I0/I3415/net049	net942	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3408/T3	I0/I3408/net049	net941	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3431/T3	I0/I3431/net049	net940	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3428/T3	I0/I3428/net049	net939	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3406/T3	I0/I3406/net049	net938	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3451/T2	BL17	net946	I0/I3451/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3441/T2	BL17	net945	I0/I3441/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3467/T2	BL17	net944	I0/I3467/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3461/T2	BL17	net943	I0/I3461/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3447/T2	BL17	net942	I0/I3447/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3440/T2	BL17	net941	I0/I3440/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3463/T2	BL17	net940	I0/I3463/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3460/T2	BL17	net939	I0/I3460/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3438/T2	BL17	net938	I0/I3438/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3759/T3	I0/I3759/net049	net937	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3759/T4	vss	I0/I3759/net13	I0/I3759/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3759/T5	I0/I3759/net13	I0/I3759/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3759/T2	BL27	net937	I0/I3759/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3727/T3	I0/I3727/net049	net937	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3727/T4	vss	I0/I3727/net13	I0/I3727/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3727/T5	I0/I3727/net13	I0/I3727/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3567/T4	vss	I0/I3567/net13	I0/I3567/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3567/T5	I0/I3567/net13	I0/I3567/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3567/T2	BL21	net937	I0/I3567/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3535/T3	I0/I3535/net049	net937	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3535/T4	vss	I0/I3535/net13	I0/I3535/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3535/T5	I0/I3535/net13	I0/I3535/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3535/T2	BL20	net937	I0/I3535/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3567/T3	I0/I3567/net049	net937	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3631/T4	vss	I0/I3631/net13	I0/I3631/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3631/T5	I0/I3631/net13	I0/I3631/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3631/T2	BL23	net937	I0/I3631/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3599/T3	I0/I3599/net049	net937	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3599/T4	vss	I0/I3599/net13	I0/I3599/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3599/T5	I0/I3599/net13	I0/I3599/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3599/T2	BL22	net937	I0/I3599/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3439/T2	BL17	net937	I0/I3439/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3407/T3	I0/I3407/net049	net937	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3407/T4	vss	I0/I3407/net13	I0/I3407/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3407/T5	I0/I3407/net13	I0/I3407/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3407/T2	BL16	net937	I0/I3407/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3631/T3	I0/I3631/net049	net937	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3766/T3	I0/I3766/net049	net936	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3766/T4	vss	I0/I3766/net13	I0/I3766/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3766/T5	I0/I3766/net13	I0/I3766/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3766/T2	BL27	net936	I0/I3766/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3734/T3	I0/I3734/net049	net936	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3734/T4	vss	I0/I3734/net13	I0/I3734/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3734/T5	I0/I3734/net13	I0/I3734/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3574/T4	vss	I0/I3574/net13	I0/I3574/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3574/T5	I0/I3574/net13	I0/I3574/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3574/T2	BL21	net936	I0/I3574/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3542/T3	I0/I3542/net049	net936	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3542/T4	vss	I0/I3542/net13	I0/I3542/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3542/T5	I0/I3542/net13	I0/I3542/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3542/T2	BL20	net936	I0/I3542/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3574/T3	I0/I3574/net049	net936	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3638/T4	vss	I0/I3638/net13	I0/I3638/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3638/T5	I0/I3638/net13	I0/I3638/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3638/T2	BL23	net936	I0/I3638/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3606/T3	I0/I3606/net049	net936	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3606/T4	vss	I0/I3606/net13	I0/I3606/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3606/T5	I0/I3606/net13	I0/I3606/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3606/T2	BL22	net936	I0/I3606/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3446/T2	BL17	net936	I0/I3446/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3414/T3	I0/I3414/net049	net936	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3414/T4	vss	I0/I3414/net13	I0/I3414/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3414/T5	I0/I3414/net13	I0/I3414/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3414/T2	BL16	net936	I0/I3414/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3638/T3	I0/I3638/net049	net936	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3768/T3	I0/I3768/net049	net935	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3768/T4	vss	I0/I3768/net13	I0/I3768/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3768/T5	I0/I3768/net13	I0/I3768/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3768/T2	BL27	net935	I0/I3768/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3736/T3	I0/I3736/net049	net935	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3736/T4	vss	I0/I3736/net13	I0/I3736/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3736/T5	I0/I3736/net13	I0/I3736/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3576/T4	vss	I0/I3576/net13	I0/I3576/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3576/T5	I0/I3576/net13	I0/I3576/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3576/T2	BL21	net935	I0/I3576/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3544/T3	I0/I3544/net049	net935	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3544/T4	vss	I0/I3544/net13	I0/I3544/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3544/T5	I0/I3544/net13	I0/I3544/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3544/T2	BL20	net935	I0/I3544/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3576/T3	I0/I3576/net049	net935	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3640/T4	vss	I0/I3640/net13	I0/I3640/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3640/T5	I0/I3640/net13	I0/I3640/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3640/T2	BL23	net935	I0/I3640/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3608/T3	I0/I3608/net049	net935	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3608/T4	vss	I0/I3608/net13	I0/I3608/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3608/T5	I0/I3608/net13	I0/I3608/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3608/T2	BL22	net935	I0/I3608/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3448/T2	BL17	net935	I0/I3448/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3416/T3	I0/I3416/net049	net935	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3416/T4	vss	I0/I3416/net13	I0/I3416/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3416/T5	I0/I3416/net13	I0/I3416/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3416/T2	BL16	net935	I0/I3416/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3640/T3	I0/I3640/net049	net935	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3774/T3	I0/I3774/net049	net934	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3774/T4	vss	I0/I3774/net13	I0/I3774/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3774/T5	I0/I3774/net13	I0/I3774/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3774/T2	BL27	net934	I0/I3774/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3742/T3	I0/I3742/net049	net934	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3742/T4	vss	I0/I3742/net13	I0/I3742/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3742/T5	I0/I3742/net13	I0/I3742/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3582/T4	vss	I0/I3582/net13	I0/I3582/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3582/T5	I0/I3582/net13	I0/I3582/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3582/T2	BL21	net934	I0/I3582/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3550/T3	I0/I3550/net049	net934	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3550/T4	vss	I0/I3550/net13	I0/I3550/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3550/T5	I0/I3550/net13	I0/I3550/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3550/T2	BL20	net934	I0/I3550/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3582/T3	I0/I3582/net049	net934	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3646/T4	vss	I0/I3646/net13	I0/I3646/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3646/T5	I0/I3646/net13	I0/I3646/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3646/T2	BL23	net934	I0/I3646/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3614/T3	I0/I3614/net049	net934	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3614/T4	vss	I0/I3614/net13	I0/I3614/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3614/T5	I0/I3614/net13	I0/I3614/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3614/T2	BL22	net934	I0/I3614/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3454/T2	BL17	net934	I0/I3454/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3422/T3	I0/I3422/net049	net934	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3422/T4	vss	I0/I3422/net13	I0/I3422/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3422/T5	I0/I3422/net13	I0/I3422/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3422/T2	BL16	net934	I0/I3422/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3646/T3	I0/I3646/net049	net934	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3776/T3	I0/I3776/net049	net933	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3776/T4	vss	I0/I3776/net13	I0/I3776/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3776/T5	I0/I3776/net13	I0/I3776/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3776/T2	BL27	net933	I0/I3776/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3744/T3	I0/I3744/net049	net933	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3744/T4	vss	I0/I3744/net13	I0/I3744/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3744/T5	I0/I3744/net13	I0/I3744/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3584/T4	vss	I0/I3584/net13	I0/I3584/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3584/T5	I0/I3584/net13	I0/I3584/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3584/T2	BL21	net933	I0/I3584/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3552/T3	I0/I3552/net049	net933	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3552/T4	vss	I0/I3552/net13	I0/I3552/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3552/T5	I0/I3552/net13	I0/I3552/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3552/T2	BL20	net933	I0/I3552/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3584/T3	I0/I3584/net049	net933	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3648/T4	vss	I0/I3648/net13	I0/I3648/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3648/T5	I0/I3648/net13	I0/I3648/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3648/T2	BL23	net933	I0/I3648/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3616/T3	I0/I3616/net049	net933	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3616/T4	vss	I0/I3616/net13	I0/I3616/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3616/T5	I0/I3616/net13	I0/I3616/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3616/T2	BL22	net933	I0/I3616/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3456/T2	BL17	net933	I0/I3456/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3424/T3	I0/I3424/net049	net933	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3424/T4	vss	I0/I3424/net13	I0/I3424/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3424/T5	I0/I3424/net13	I0/I3424/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3424/T2	BL16	net933	I0/I3424/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3648/T3	I0/I3648/net049	net933	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3765/T3	I0/I3765/net049	net932	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3765/T4	vss	I0/I3765/net13	I0/I3765/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3765/T5	I0/I3765/net13	I0/I3765/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3765/T2	BL27	net932	I0/I3765/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3733/T3	I0/I3733/net049	net932	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3733/T4	vss	I0/I3733/net13	I0/I3733/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3733/T5	I0/I3733/net13	I0/I3733/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3573/T4	vss	I0/I3573/net13	I0/I3573/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3573/T5	I0/I3573/net13	I0/I3573/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3573/T2	BL21	net932	I0/I3573/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3541/T3	I0/I3541/net049	net932	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3541/T4	vss	I0/I3541/net13	I0/I3541/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3541/T5	I0/I3541/net13	I0/I3541/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3541/T2	BL20	net932	I0/I3541/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3573/T3	I0/I3573/net049	net932	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3637/T4	vss	I0/I3637/net13	I0/I3637/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3637/T5	I0/I3637/net13	I0/I3637/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3637/T2	BL23	net932	I0/I3637/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3605/T3	I0/I3605/net049	net932	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3605/T4	vss	I0/I3605/net13	I0/I3605/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3605/T5	I0/I3605/net13	I0/I3605/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3605/T2	BL22	net932	I0/I3605/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3445/T2	BL17	net932	I0/I3445/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3413/T3	I0/I3413/net049	net932	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3413/T4	vss	I0/I3413/net13	I0/I3413/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3413/T5	I0/I3413/net13	I0/I3413/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3413/T2	BL16	net932	I0/I3413/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3637/T3	I0/I3637/net049	net932	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3779/T3	I0/I3779/net049	net931	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3779/T4	vss	I0/I3779/net13	I0/I3779/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3779/T5	I0/I3779/net13	I0/I3779/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3779/T2	BL27	net931	I0/I3779/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3747/T3	I0/I3747/net049	net931	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3747/T4	vss	I0/I3747/net13	I0/I3747/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3747/T5	I0/I3747/net13	I0/I3747/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3587/T4	vss	I0/I3587/net13	I0/I3587/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3587/T5	I0/I3587/net13	I0/I3587/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3587/T2	BL21	net931	I0/I3587/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3555/T3	I0/I3555/net049	net931	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3555/T4	vss	I0/I3555/net13	I0/I3555/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3555/T5	I0/I3555/net13	I0/I3555/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3555/T2	BL20	net931	I0/I3555/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3587/T3	I0/I3587/net049	net931	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3651/T4	vss	I0/I3651/net13	I0/I3651/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3651/T5	I0/I3651/net13	I0/I3651/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3651/T2	BL23	net931	I0/I3651/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3619/T3	I0/I3619/net049	net931	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3619/T4	vss	I0/I3619/net13	I0/I3619/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3619/T5	I0/I3619/net13	I0/I3619/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3619/T2	BL22	net931	I0/I3619/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3459/T2	BL17	net931	I0/I3459/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3427/T3	I0/I3427/net049	net931	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3427/T4	vss	I0/I3427/net13	I0/I3427/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3427/T5	I0/I3427/net13	I0/I3427/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3427/T2	BL16	net931	I0/I3427/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3651/T3	I0/I3651/net049	net931	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3773/T3	I0/I3773/net049	net930	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3773/T4	vss	I0/I3773/net13	I0/I3773/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3773/T5	I0/I3773/net13	I0/I3773/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3773/T2	BL27	net930	I0/I3773/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3741/T3	I0/I3741/net049	net930	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3741/T4	vss	I0/I3741/net13	I0/I3741/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3741/T5	I0/I3741/net13	I0/I3741/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3581/T4	vss	I0/I3581/net13	I0/I3581/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3581/T5	I0/I3581/net13	I0/I3581/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3581/T2	BL21	net930	I0/I3581/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3549/T3	I0/I3549/net049	net930	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3549/T4	vss	I0/I3549/net13	I0/I3549/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3549/T5	I0/I3549/net13	I0/I3549/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3549/T2	BL20	net930	I0/I3549/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3581/T3	I0/I3581/net049	net930	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3645/T4	vss	I0/I3645/net13	I0/I3645/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3645/T5	I0/I3645/net13	I0/I3645/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3645/T2	BL23	net930	I0/I3645/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3613/T3	I0/I3613/net049	net930	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3613/T4	vss	I0/I3613/net13	I0/I3613/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3613/T5	I0/I3613/net13	I0/I3613/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3613/T2	BL22	net930	I0/I3613/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3453/T2	BL17	net930	I0/I3453/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3421/T3	I0/I3421/net049	net930	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3421/T4	vss	I0/I3421/net13	I0/I3421/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3421/T5	I0/I3421/net13	I0/I3421/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3421/T2	BL16	net930	I0/I3421/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3645/T3	I0/I3645/net049	net930	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3777/T3	I0/I3777/net049	net929	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3777/T4	vss	I0/I3777/net13	I0/I3777/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3777/T5	I0/I3777/net13	I0/I3777/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3777/T2	BL27	net929	I0/I3777/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3745/T3	I0/I3745/net049	net929	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3745/T4	vss	I0/I3745/net13	I0/I3745/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3745/T5	I0/I3745/net13	I0/I3745/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3585/T4	vss	I0/I3585/net13	I0/I3585/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3585/T5	I0/I3585/net13	I0/I3585/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3585/T2	BL21	net929	I0/I3585/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3553/T3	I0/I3553/net049	net929	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3553/T4	vss	I0/I3553/net13	I0/I3553/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3553/T5	I0/I3553/net13	I0/I3553/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3553/T2	BL20	net929	I0/I3553/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3585/T3	I0/I3585/net049	net929	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3649/T4	vss	I0/I3649/net13	I0/I3649/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3649/T5	I0/I3649/net13	I0/I3649/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3649/T2	BL23	net929	I0/I3649/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3617/T3	I0/I3617/net049	net929	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3617/T4	vss	I0/I3617/net13	I0/I3617/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3617/T5	I0/I3617/net13	I0/I3617/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3617/T2	BL22	net929	I0/I3617/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3457/T2	BL17	net929	I0/I3457/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3425/T3	I0/I3425/net049	net929	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3425/T4	vss	I0/I3425/net13	I0/I3425/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3425/T5	I0/I3425/net13	I0/I3425/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3425/T2	BL16	net929	I0/I3425/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3649/T3	I0/I3649/net049	net929	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3789/T3	I0/I3789/net049	net928	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3789/T4	vss	I0/I3789/net13	I0/I3789/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3789/T5	I0/I3789/net13	I0/I3789/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3789/T2	BL27	net928	I0/I3789/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3757/T3	I0/I3757/net049	net928	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3757/T4	vss	I0/I3757/net13	I0/I3757/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3757/T5	I0/I3757/net13	I0/I3757/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3597/T4	vss	I0/I3597/net13	I0/I3597/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3597/T5	I0/I3597/net13	I0/I3597/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3597/T2	BL21	net928	I0/I3597/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3565/T3	I0/I3565/net049	net928	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3565/T4	vss	I0/I3565/net13	I0/I3565/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3565/T5	I0/I3565/net13	I0/I3565/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3565/T2	BL20	net928	I0/I3565/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3597/T3	I0/I3597/net049	net928	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3661/T4	vss	I0/I3661/net13	I0/I3661/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3661/T5	I0/I3661/net13	I0/I3661/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3661/T2	BL23	net928	I0/I3661/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3629/T3	I0/I3629/net049	net928	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3629/T4	vss	I0/I3629/net13	I0/I3629/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3629/T5	I0/I3629/net13	I0/I3629/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3629/T2	BL22	net928	I0/I3629/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3469/T2	BL17	net928	I0/I3469/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3437/T3	I0/I3437/net049	net928	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3437/T4	vss	I0/I3437/net13	I0/I3437/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3437/T5	I0/I3437/net13	I0/I3437/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3437/T2	BL16	net928	I0/I3437/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3661/T3	I0/I3661/net049	net928	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3775/T3	I0/I3775/net049	net927	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3775/T4	vss	I0/I3775/net13	I0/I3775/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3775/T5	I0/I3775/net13	I0/I3775/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3775/T2	BL27	net927	I0/I3775/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3743/T3	I0/I3743/net049	net927	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3743/T4	vss	I0/I3743/net13	I0/I3743/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3743/T5	I0/I3743/net13	I0/I3743/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3583/T4	vss	I0/I3583/net13	I0/I3583/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3583/T5	I0/I3583/net13	I0/I3583/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3583/T2	BL21	net927	I0/I3583/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3551/T3	I0/I3551/net049	net927	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3551/T4	vss	I0/I3551/net13	I0/I3551/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3551/T5	I0/I3551/net13	I0/I3551/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3551/T2	BL20	net927	I0/I3551/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3583/T3	I0/I3583/net049	net927	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3647/T4	vss	I0/I3647/net13	I0/I3647/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3647/T5	I0/I3647/net13	I0/I3647/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3647/T2	BL23	net927	I0/I3647/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3615/T3	I0/I3615/net049	net927	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3615/T4	vss	I0/I3615/net13	I0/I3615/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3615/T5	I0/I3615/net13	I0/I3615/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3615/T2	BL22	net927	I0/I3615/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3455/T2	BL17	net927	I0/I3455/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3423/T3	I0/I3423/net049	net927	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3423/T4	vss	I0/I3423/net13	I0/I3423/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3423/T5	I0/I3423/net13	I0/I3423/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3423/T2	BL16	net927	I0/I3423/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3647/T3	I0/I3647/net049	net927	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3786/T3	I0/I3786/net049	net926	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3786/T4	vss	I0/I3786/net13	I0/I3786/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3786/T5	I0/I3786/net13	I0/I3786/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3786/T2	BL27	net926	I0/I3786/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3754/T3	I0/I3754/net049	net926	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3754/T4	vss	I0/I3754/net13	I0/I3754/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3754/T5	I0/I3754/net13	I0/I3754/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3594/T4	vss	I0/I3594/net13	I0/I3594/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3594/T5	I0/I3594/net13	I0/I3594/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3594/T2	BL21	net926	I0/I3594/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3562/T3	I0/I3562/net049	net926	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3562/T4	vss	I0/I3562/net13	I0/I3562/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3562/T5	I0/I3562/net13	I0/I3562/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3562/T2	BL20	net926	I0/I3562/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3594/T3	I0/I3594/net049	net926	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3658/T4	vss	I0/I3658/net13	I0/I3658/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3658/T5	I0/I3658/net13	I0/I3658/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3658/T2	BL23	net926	I0/I3658/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3626/T3	I0/I3626/net049	net926	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3626/T4	vss	I0/I3626/net13	I0/I3626/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3626/T5	I0/I3626/net13	I0/I3626/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3626/T2	BL22	net926	I0/I3626/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3466/T2	BL17	net926	I0/I3466/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3434/T3	I0/I3434/net049	net926	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3434/T4	vss	I0/I3434/net13	I0/I3434/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3434/T5	I0/I3434/net13	I0/I3434/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3434/T2	BL16	net926	I0/I3434/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3658/T3	I0/I3658/net049	net926	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3785/T3	I0/I3785/net049	net925	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3785/T4	vss	I0/I3785/net13	I0/I3785/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3785/T5	I0/I3785/net13	I0/I3785/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3785/T2	BL27	net925	I0/I3785/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3753/T3	I0/I3753/net049	net925	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3753/T4	vss	I0/I3753/net13	I0/I3753/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3753/T5	I0/I3753/net13	I0/I3753/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3593/T4	vss	I0/I3593/net13	I0/I3593/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3593/T5	I0/I3593/net13	I0/I3593/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3593/T2	BL21	net925	I0/I3593/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3561/T3	I0/I3561/net049	net925	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3561/T4	vss	I0/I3561/net13	I0/I3561/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3561/T5	I0/I3561/net13	I0/I3561/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3561/T2	BL20	net925	I0/I3561/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3593/T3	I0/I3593/net049	net925	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3657/T4	vss	I0/I3657/net13	I0/I3657/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3657/T5	I0/I3657/net13	I0/I3657/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3657/T2	BL23	net925	I0/I3657/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3625/T3	I0/I3625/net049	net925	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3625/T4	vss	I0/I3625/net13	I0/I3625/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3625/T5	I0/I3625/net13	I0/I3625/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3625/T2	BL22	net925	I0/I3625/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3465/T2	BL17	net925	I0/I3465/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3433/T3	I0/I3433/net049	net925	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3433/T4	vss	I0/I3433/net13	I0/I3433/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3433/T5	I0/I3433/net13	I0/I3433/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3433/T2	BL16	net925	I0/I3433/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3657/T3	I0/I3657/net049	net925	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3762/T3	I0/I3762/net049	net924	BL27bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3762/T4	vss	I0/I3762/net13	I0/I3762/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3762/T5	I0/I3762/net13	I0/I3762/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3762/T2	BL27	net924	I0/I3762/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3730/T3	I0/I3730/net049	net924	BL26bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3730/T4	vss	I0/I3730/net13	I0/I3730/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3730/T5	I0/I3730/net13	I0/I3730/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3570/T4	vss	I0/I3570/net13	I0/I3570/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3570/T5	I0/I3570/net13	I0/I3570/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3570/T2	BL21	net924	I0/I3570/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3538/T3	I0/I3538/net049	net924	BL20bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3538/T4	vss	I0/I3538/net13	I0/I3538/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3538/T5	I0/I3538/net13	I0/I3538/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3538/T2	BL20	net924	I0/I3538/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3570/T3	I0/I3570/net049	net924	BL21bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3634/T4	vss	I0/I3634/net13	I0/I3634/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3634/T5	I0/I3634/net13	I0/I3634/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3634/T2	BL23	net924	I0/I3634/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3602/T3	I0/I3602/net049	net924	BL22bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3602/T4	vss	I0/I3602/net13	I0/I3602/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3602/T5	I0/I3602/net13	I0/I3602/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3602/T2	BL22	net924	I0/I3602/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3442/T2	BL17	net924	I0/I3442/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3410/T3	I0/I3410/net049	net924	BL16bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3410/T4	vss	I0/I3410/net13	I0/I3410/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3410/T5	I0/I3410/net13	I0/I3410/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3410/T2	BL16	net924	I0/I3410/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3634/T3	I0/I3634/net049	net924	BL23bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI80/T1	p6bar	y2	BL21bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI81/T1	BL21	y2	p6	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI82/T1	p6bar	y1	BL20bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI83/T1	BL20	y1	p6	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI84/T1	p7bar	y4	BL27bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI85/T1	BL27	y4	p7	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI86/T1	p7bar	y3	BL26bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T2	I5/net23	p5	I5/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T3	I5/net20	p5bar	I5/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T4	vss	vdd	I5/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T8	vss	I5/net20	I5/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T7	data4	I5/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T11	I27/net23	data4	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T16	I27/net15	net680	p5	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T17	vss	I27/net23	I27/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T19	I27/net7	p5	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T18	p5bar	net680	I27/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T2	I6/net23	p6	I6/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T3	I6/net20	p6bar	I6/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T16	I26/net15	net680	p4	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI77/T1	BL23	y4	p6	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T17	vss	I26/net23	I26/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T19	I26/net7	p4	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI78/T1	p6bar	y3	BL22bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T18	p4bar	net680	I26/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI79/T1	BL22	y3	p6	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI73/T1	BL17	y2	p5	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T3	I4/net20	p4bar	I4/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI74/T1	p5bar	y1	BL16bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T4	vss	vdd	I4/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T8	vss	I4/net20	I4/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI75/T1	BL16	y1	p5	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T7	data3	I4/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI76/T1	p6bar	y4	BL23bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T11	I26/net23	data3	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T2	I4/net23	p4	I4/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3452/T3	I0/I3452/net049	net955	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3444/T3	I0/I3444/net049	net954	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3452/T4	vss	I0/I3452/net13	I0/I3452/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3444/T4	vss	I0/I3444/net13	I0/I3444/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3452/T5	I0/I3452/net13	I0/I3452/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3444/T5	I0/I3444/net13	I0/I3444/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3443/T3	I0/I3443/net049	net953	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3468/T3	I0/I3468/net049	net952	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3443/T4	vss	I0/I3443/net13	I0/I3443/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3468/T4	vss	I0/I3468/net13	I0/I3468/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3443/T5	I0/I3443/net13	I0/I3443/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3468/T5	I0/I3468/net13	I0/I3468/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3449/T3	I0/I3449/net049	net951	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3449/T4	vss	I0/I3449/net13	I0/I3449/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3449/T5	I0/I3449/net13	I0/I3449/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3464/T3	I0/I3464/net049	net950	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3462/T3	I0/I3462/net049	net949	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3464/T4	vss	I0/I3464/net13	I0/I3464/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3462/T4	vss	I0/I3462/net13	I0/I3462/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3464/T5	I0/I3464/net13	I0/I3464/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3462/T5	I0/I3462/net13	I0/I3462/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3458/T3	I0/I3458/net049	net948	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3450/T3	I0/I3450/net049	net947	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3458/T4	vss	I0/I3458/net13	I0/I3458/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3450/T4	vss	I0/I3450/net13	I0/I3450/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3458/T5	I0/I3458/net13	I0/I3458/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3450/T5	I0/I3450/net13	I0/I3450/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3484/T2	BL18	net955	I0/I3484/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3476/T2	BL18	net954	I0/I3476/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3475/T2	BL18	net953	I0/I3475/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3500/T2	BL18	net952	I0/I3500/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3481/T2	BL18	net951	I0/I3481/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3496/T2	BL18	net950	I0/I3496/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3494/T2	BL18	net949	I0/I3494/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3490/T2	BL18	net948	I0/I3490/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3482/T2	BL18	net947	I0/I3482/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3484/T5	I0/I3484/net13	I0/I3484/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3476/T5	I0/I3476/net13	I0/I3476/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3475/T5	I0/I3475/net13	I0/I3475/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3500/T5	I0/I3500/net13	I0/I3500/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3481/T5	I0/I3481/net13	I0/I3481/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3496/T5	I0/I3496/net13	I0/I3496/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3494/T5	I0/I3494/net13	I0/I3494/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3490/T5	I0/I3490/net13	I0/I3490/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3482/T5	I0/I3482/net13	I0/I3482/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3484/T4	vss	I0/I3484/net13	I0/I3484/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3476/T4	vss	I0/I3476/net13	I0/I3476/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3475/T4	vss	I0/I3475/net13	I0/I3475/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3500/T4	vss	I0/I3500/net13	I0/I3500/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3481/T4	vss	I0/I3481/net13	I0/I3481/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3496/T4	vss	I0/I3496/net13	I0/I3496/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3494/T4	vss	I0/I3494/net13	I0/I3494/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3490/T4	vss	I0/I3490/net13	I0/I3490/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3482/T4	vss	I0/I3482/net13	I0/I3482/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3484/T3	I0/I3484/net049	net955	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3476/T3	I0/I3476/net049	net954	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3475/T3	I0/I3475/net049	net953	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3500/T3	I0/I3500/net049	net952	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3481/T3	I0/I3481/net049	net951	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3496/T3	I0/I3496/net049	net950	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3494/T3	I0/I3494/net049	net949	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3490/T3	I0/I3490/net049	net948	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3482/T3	I0/I3482/net049	net947	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3516/T2	BL19	net955	I0/I3516/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3508/T2	BL19	net954	I0/I3508/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3507/T2	BL19	net953	I0/I3507/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3532/T2	BL19	net952	I0/I3532/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3513/T2	BL19	net951	I0/I3513/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3528/T2	BL19	net950	I0/I3528/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3526/T2	BL19	net949	I0/I3526/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3522/T2	BL19	net948	I0/I3522/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3514/T2	BL19	net947	I0/I3514/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3516/T5	I0/I3516/net13	I0/I3516/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3508/T5	I0/I3508/net13	I0/I3508/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3507/T5	I0/I3507/net13	I0/I3507/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3532/T5	I0/I3532/net13	I0/I3532/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3513/T5	I0/I3513/net13	I0/I3513/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3528/T5	I0/I3528/net13	I0/I3528/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3526/T5	I0/I3526/net13	I0/I3526/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3522/T5	I0/I3522/net13	I0/I3522/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3514/T5	I0/I3514/net13	I0/I3514/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3516/T4	vss	I0/I3516/net13	I0/I3516/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3508/T4	vss	I0/I3508/net13	I0/I3508/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3507/T4	vss	I0/I3507/net13	I0/I3507/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3532/T4	vss	I0/I3532/net13	I0/I3532/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3513/T4	vss	I0/I3513/net13	I0/I3513/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3528/T4	vss	I0/I3528/net13	I0/I3528/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3526/T4	vss	I0/I3526/net13	I0/I3526/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3522/T4	vss	I0/I3522/net13	I0/I3522/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3514/T4	vss	I0/I3514/net13	I0/I3514/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3516/T3	I0/I3516/net049	net955	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3508/T3	I0/I3508/net049	net954	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3507/T3	I0/I3507/net049	net953	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3532/T3	I0/I3532/net049	net952	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3513/T3	I0/I3513/net049	net951	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3528/T3	I0/I3528/net049	net950	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3526/T3	I0/I3526/net049	net949	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3522/T3	I0/I3522/net049	net948	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3514/T3	I0/I3514/net049	net947	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3292/T4	vss	I0/I3292/net13	I0/I3292/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3284/T4	vss	I0/I3284/net13	I0/I3284/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3292/T5	I0/I3292/net13	I0/I3292/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3284/T5	I0/I3284/net13	I0/I3284/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3292/T2	BL12	net955	I0/I3292/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3284/T2	BL12	net954	I0/I3284/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3283/T4	vss	I0/I3283/net13	I0/I3283/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3308/T4	vss	I0/I3308/net13	I0/I3308/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3283/T5	I0/I3283/net13	I0/I3283/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3308/T5	I0/I3308/net13	I0/I3308/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3283/T2	BL12	net953	I0/I3283/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3308/T2	BL12	net952	I0/I3308/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3289/T4	vss	I0/I3289/net13	I0/I3289/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3289/T5	I0/I3289/net13	I0/I3289/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3289/T2	BL12	net951	I0/I3289/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3304/T4	vss	I0/I3304/net13	I0/I3304/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3302/T4	vss	I0/I3302/net13	I0/I3302/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3304/T5	I0/I3304/net13	I0/I3304/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3302/T5	I0/I3302/net13	I0/I3302/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3304/T2	BL12	net950	I0/I3304/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3302/T2	BL12	net949	I0/I3302/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3298/T4	vss	I0/I3298/net13	I0/I3298/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3290/T4	vss	I0/I3290/net13	I0/I3290/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3298/T5	I0/I3298/net13	I0/I3298/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3290/T5	I0/I3290/net13	I0/I3290/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3298/T2	BL12	net948	I0/I3298/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3290/T2	BL12	net947	I0/I3290/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3292/T3	I0/I3292/net049	net955	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3284/T3	I0/I3284/net049	net954	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3283/T3	I0/I3283/net049	net953	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3308/T3	I0/I3308/net049	net952	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3289/T3	I0/I3289/net049	net951	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3304/T3	I0/I3304/net049	net950	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3302/T3	I0/I3302/net049	net949	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3298/T3	I0/I3298/net049	net948	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3290/T3	I0/I3290/net049	net947	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3324/T2	BL13	net955	I0/I3324/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3316/T2	BL13	net954	I0/I3316/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3315/T2	BL13	net953	I0/I3315/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3340/T2	BL13	net952	I0/I3340/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3321/T2	BL13	net951	I0/I3321/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3336/T2	BL13	net950	I0/I3336/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3334/T2	BL13	net949	I0/I3334/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3330/T2	BL13	net948	I0/I3330/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3322/T2	BL13	net947	I0/I3322/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3324/T5	I0/I3324/net13	I0/I3324/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3316/T5	I0/I3316/net13	I0/I3316/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3315/T5	I0/I3315/net13	I0/I3315/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3340/T5	I0/I3340/net13	I0/I3340/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3321/T5	I0/I3321/net13	I0/I3321/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3336/T5	I0/I3336/net13	I0/I3336/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3334/T5	I0/I3334/net13	I0/I3334/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3330/T5	I0/I3330/net13	I0/I3330/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3322/T5	I0/I3322/net13	I0/I3322/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3324/T4	vss	I0/I3324/net13	I0/I3324/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3316/T4	vss	I0/I3316/net13	I0/I3316/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3315/T4	vss	I0/I3315/net13	I0/I3315/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3340/T4	vss	I0/I3340/net13	I0/I3340/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3321/T4	vss	I0/I3321/net13	I0/I3321/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3336/T4	vss	I0/I3336/net13	I0/I3336/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3334/T4	vss	I0/I3334/net13	I0/I3334/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3330/T4	vss	I0/I3330/net13	I0/I3330/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3322/T4	vss	I0/I3322/net13	I0/I3322/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3324/T3	I0/I3324/net049	net955	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3316/T3	I0/I3316/net049	net954	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3315/T3	I0/I3315/net049	net953	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3340/T3	I0/I3340/net049	net952	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3321/T3	I0/I3321/net049	net951	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3336/T3	I0/I3336/net049	net950	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3334/T3	I0/I3334/net049	net949	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3330/T3	I0/I3330/net049	net948	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3322/T3	I0/I3322/net049	net947	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3356/T4	vss	I0/I3356/net13	I0/I3356/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3348/T4	vss	I0/I3348/net13	I0/I3348/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3356/T5	I0/I3356/net13	I0/I3356/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3348/T5	I0/I3348/net13	I0/I3348/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3356/T2	BL14	net955	I0/I3356/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3348/T2	BL14	net954	I0/I3348/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3347/T4	vss	I0/I3347/net13	I0/I3347/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3372/T4	vss	I0/I3372/net13	I0/I3372/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3347/T5	I0/I3347/net13	I0/I3347/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3372/T5	I0/I3372/net13	I0/I3372/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3347/T2	BL14	net953	I0/I3347/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3372/T2	BL14	net952	I0/I3372/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3353/T4	vss	I0/I3353/net13	I0/I3353/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3353/T5	I0/I3353/net13	I0/I3353/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3353/T2	BL14	net951	I0/I3353/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3368/T4	vss	I0/I3368/net13	I0/I3368/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3366/T4	vss	I0/I3366/net13	I0/I3366/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3368/T5	I0/I3368/net13	I0/I3368/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3366/T5	I0/I3366/net13	I0/I3366/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3368/T2	BL14	net950	I0/I3368/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3366/T2	BL14	net949	I0/I3366/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3362/T4	vss	I0/I3362/net13	I0/I3362/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3354/T4	vss	I0/I3354/net13	I0/I3354/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3362/T5	I0/I3362/net13	I0/I3362/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3354/T5	I0/I3354/net13	I0/I3354/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3362/T2	BL14	net948	I0/I3362/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3354/T2	BL14	net947	I0/I3354/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3356/T3	I0/I3356/net049	net955	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3348/T3	I0/I3348/net049	net954	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3347/T3	I0/I3347/net049	net953	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3372/T3	I0/I3372/net049	net952	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3353/T3	I0/I3353/net049	net951	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3368/T3	I0/I3368/net049	net950	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3366/T3	I0/I3366/net049	net949	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3362/T3	I0/I3362/net049	net948	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3354/T3	I0/I3354/net049	net947	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3388/T2	BL15	net955	I0/I3388/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3380/T2	BL15	net954	I0/I3380/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3379/T2	BL15	net953	I0/I3379/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3404/T2	BL15	net952	I0/I3404/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3385/T2	BL15	net951	I0/I3385/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3400/T2	BL15	net950	I0/I3400/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3398/T2	BL15	net949	I0/I3398/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3394/T2	BL15	net948	I0/I3394/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3386/T2	BL15	net947	I0/I3386/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3388/T5	I0/I3388/net13	I0/I3388/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3380/T5	I0/I3380/net13	I0/I3380/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3379/T5	I0/I3379/net13	I0/I3379/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3404/T5	I0/I3404/net13	I0/I3404/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3385/T5	I0/I3385/net13	I0/I3385/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3400/T5	I0/I3400/net13	I0/I3400/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3398/T5	I0/I3398/net13	I0/I3398/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3394/T5	I0/I3394/net13	I0/I3394/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3386/T5	I0/I3386/net13	I0/I3386/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3388/T4	vss	I0/I3388/net13	I0/I3388/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3380/T4	vss	I0/I3380/net13	I0/I3380/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3379/T4	vss	I0/I3379/net13	I0/I3379/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3404/T4	vss	I0/I3404/net13	I0/I3404/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3385/T4	vss	I0/I3385/net13	I0/I3385/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3400/T4	vss	I0/I3400/net13	I0/I3400/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3398/T4	vss	I0/I3398/net13	I0/I3398/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3394/T4	vss	I0/I3394/net13	I0/I3394/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3386/T4	vss	I0/I3386/net13	I0/I3386/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3388/T3	I0/I3388/net049	net955	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3380/T3	I0/I3380/net049	net954	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3379/T3	I0/I3379/net049	net953	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3404/T3	I0/I3404/net049	net952	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3385/T3	I0/I3385/net049	net951	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3400/T3	I0/I3400/net049	net950	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3398/T3	I0/I3398/net049	net949	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3394/T3	I0/I3394/net049	net948	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3386/T3	I0/I3386/net049	net947	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3100/T2	BL8	net955	I0/I3100/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3092/T2	BL8	net954	I0/I3092/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3091/T2	BL8	net953	I0/I3091/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3116/T2	BL8	net952	I0/I3116/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3097/T2	BL8	net951	I0/I3097/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3112/T2	BL8	net950	I0/I3112/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3110/T2	BL8	net949	I0/I3110/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3106/T2	BL8	net948	I0/I3106/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3098/T2	BL8	net947	I0/I3098/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3451/T3	I0/I3451/net049	net946	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3441/T3	I0/I3441/net049	net945	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3451/T4	vss	I0/I3451/net13	I0/I3451/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3441/T4	vss	I0/I3441/net13	I0/I3441/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3451/T5	I0/I3451/net13	I0/I3451/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3441/T5	I0/I3441/net13	I0/I3441/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3467/T3	I0/I3467/net049	net944	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3461/T3	I0/I3461/net049	net943	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3467/T4	vss	I0/I3467/net13	I0/I3467/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3461/T4	vss	I0/I3461/net13	I0/I3461/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3467/T5	I0/I3467/net13	I0/I3467/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3461/T5	I0/I3461/net13	I0/I3461/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3447/T3	I0/I3447/net049	net942	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3447/T4	vss	I0/I3447/net13	I0/I3447/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3447/T5	I0/I3447/net13	I0/I3447/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3440/T3	I0/I3440/net049	net941	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3463/T3	I0/I3463/net049	net940	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3440/T4	vss	I0/I3440/net13	I0/I3440/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3463/T4	vss	I0/I3463/net13	I0/I3463/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3440/T5	I0/I3440/net13	I0/I3440/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3463/T5	I0/I3463/net13	I0/I3463/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3460/T3	I0/I3460/net049	net939	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3438/T3	I0/I3438/net049	net938	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3460/T4	vss	I0/I3460/net13	I0/I3460/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3438/T4	vss	I0/I3438/net13	I0/I3438/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3460/T5	I0/I3460/net13	I0/I3460/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3438/T5	I0/I3438/net13	I0/I3438/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3483/T2	BL18	net946	I0/I3483/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3473/T2	BL18	net945	I0/I3473/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3499/T2	BL18	net944	I0/I3499/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3493/T2	BL18	net943	I0/I3493/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3479/T2	BL18	net942	I0/I3479/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3472/T2	BL18	net941	I0/I3472/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3495/T2	BL18	net940	I0/I3495/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3492/T2	BL18	net939	I0/I3492/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3470/T2	BL18	net938	I0/I3470/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3483/T5	I0/I3483/net13	I0/I3483/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3473/T5	I0/I3473/net13	I0/I3473/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3499/T5	I0/I3499/net13	I0/I3499/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3493/T5	I0/I3493/net13	I0/I3493/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3479/T5	I0/I3479/net13	I0/I3479/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3472/T5	I0/I3472/net13	I0/I3472/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3495/T5	I0/I3495/net13	I0/I3495/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3492/T5	I0/I3492/net13	I0/I3492/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3470/T5	I0/I3470/net13	I0/I3470/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3483/T4	vss	I0/I3483/net13	I0/I3483/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3473/T4	vss	I0/I3473/net13	I0/I3473/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3499/T4	vss	I0/I3499/net13	I0/I3499/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3493/T4	vss	I0/I3493/net13	I0/I3493/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3479/T4	vss	I0/I3479/net13	I0/I3479/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3472/T4	vss	I0/I3472/net13	I0/I3472/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3495/T4	vss	I0/I3495/net13	I0/I3495/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3492/T4	vss	I0/I3492/net13	I0/I3492/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3470/T4	vss	I0/I3470/net13	I0/I3470/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3483/T3	I0/I3483/net049	net946	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3473/T3	I0/I3473/net049	net945	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3499/T3	I0/I3499/net049	net944	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3493/T3	I0/I3493/net049	net943	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3479/T3	I0/I3479/net049	net942	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3472/T3	I0/I3472/net049	net941	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3495/T3	I0/I3495/net049	net940	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3492/T3	I0/I3492/net049	net939	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3470/T3	I0/I3470/net049	net938	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3515/T2	BL19	net946	I0/I3515/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3505/T2	BL19	net945	I0/I3505/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3531/T2	BL19	net944	I0/I3531/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3525/T2	BL19	net943	I0/I3525/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3511/T2	BL19	net942	I0/I3511/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3504/T2	BL19	net941	I0/I3504/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3527/T2	BL19	net940	I0/I3527/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3524/T2	BL19	net939	I0/I3524/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3502/T2	BL19	net938	I0/I3502/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3515/T5	I0/I3515/net13	I0/I3515/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3505/T5	I0/I3505/net13	I0/I3505/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3531/T5	I0/I3531/net13	I0/I3531/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3525/T5	I0/I3525/net13	I0/I3525/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3511/T5	I0/I3511/net13	I0/I3511/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3504/T5	I0/I3504/net13	I0/I3504/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3527/T5	I0/I3527/net13	I0/I3527/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3524/T5	I0/I3524/net13	I0/I3524/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3502/T5	I0/I3502/net13	I0/I3502/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3515/T4	vss	I0/I3515/net13	I0/I3515/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3505/T4	vss	I0/I3505/net13	I0/I3505/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3531/T4	vss	I0/I3531/net13	I0/I3531/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3525/T4	vss	I0/I3525/net13	I0/I3525/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3511/T4	vss	I0/I3511/net13	I0/I3511/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3504/T4	vss	I0/I3504/net13	I0/I3504/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3527/T4	vss	I0/I3527/net13	I0/I3527/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3524/T4	vss	I0/I3524/net13	I0/I3524/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3502/T4	vss	I0/I3502/net13	I0/I3502/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3515/T3	I0/I3515/net049	net946	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3505/T3	I0/I3505/net049	net945	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3531/T3	I0/I3531/net049	net944	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3525/T3	I0/I3525/net049	net943	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3511/T3	I0/I3511/net049	net942	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3504/T3	I0/I3504/net049	net941	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3527/T3	I0/I3527/net049	net940	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3524/T3	I0/I3524/net049	net939	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3502/T3	I0/I3502/net049	net938	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3291/T4	vss	I0/I3291/net13	I0/I3291/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3281/T4	vss	I0/I3281/net13	I0/I3281/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3291/T5	I0/I3291/net13	I0/I3291/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3281/T5	I0/I3281/net13	I0/I3281/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3291/T2	BL12	net946	I0/I3291/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3281/T2	BL12	net945	I0/I3281/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3307/T4	vss	I0/I3307/net13	I0/I3307/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3301/T4	vss	I0/I3301/net13	I0/I3301/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3307/T5	I0/I3307/net13	I0/I3307/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3301/T5	I0/I3301/net13	I0/I3301/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3307/T2	BL12	net944	I0/I3307/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3301/T2	BL12	net943	I0/I3301/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3287/T4	vss	I0/I3287/net13	I0/I3287/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3287/T5	I0/I3287/net13	I0/I3287/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3287/T2	BL12	net942	I0/I3287/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3280/T4	vss	I0/I3280/net13	I0/I3280/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3303/T4	vss	I0/I3303/net13	I0/I3303/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3280/T5	I0/I3280/net13	I0/I3280/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3303/T5	I0/I3303/net13	I0/I3303/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3280/T2	BL12	net941	I0/I3280/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3303/T2	BL12	net940	I0/I3303/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3300/T4	vss	I0/I3300/net13	I0/I3300/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3278/T4	vss	I0/I3278/net13	I0/I3278/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3300/T5	I0/I3300/net13	I0/I3300/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3278/T5	I0/I3278/net13	I0/I3278/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3300/T2	BL12	net939	I0/I3300/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3278/T2	BL12	net938	I0/I3278/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3291/T3	I0/I3291/net049	net946	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3281/T3	I0/I3281/net049	net945	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3307/T3	I0/I3307/net049	net944	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3301/T3	I0/I3301/net049	net943	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3287/T3	I0/I3287/net049	net942	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3280/T3	I0/I3280/net049	net941	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3303/T3	I0/I3303/net049	net940	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3300/T3	I0/I3300/net049	net939	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3278/T3	I0/I3278/net049	net938	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3323/T2	BL13	net946	I0/I3323/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3313/T2	BL13	net945	I0/I3313/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3339/T2	BL13	net944	I0/I3339/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3333/T2	BL13	net943	I0/I3333/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3319/T2	BL13	net942	I0/I3319/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3312/T2	BL13	net941	I0/I3312/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3335/T2	BL13	net940	I0/I3335/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3332/T2	BL13	net939	I0/I3332/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3310/T2	BL13	net938	I0/I3310/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3323/T5	I0/I3323/net13	I0/I3323/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3313/T5	I0/I3313/net13	I0/I3313/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3339/T5	I0/I3339/net13	I0/I3339/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3333/T5	I0/I3333/net13	I0/I3333/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3319/T5	I0/I3319/net13	I0/I3319/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3312/T5	I0/I3312/net13	I0/I3312/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3335/T5	I0/I3335/net13	I0/I3335/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3332/T5	I0/I3332/net13	I0/I3332/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3310/T5	I0/I3310/net13	I0/I3310/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3323/T4	vss	I0/I3323/net13	I0/I3323/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3313/T4	vss	I0/I3313/net13	I0/I3313/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3339/T4	vss	I0/I3339/net13	I0/I3339/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3333/T4	vss	I0/I3333/net13	I0/I3333/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3319/T4	vss	I0/I3319/net13	I0/I3319/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3312/T4	vss	I0/I3312/net13	I0/I3312/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3335/T4	vss	I0/I3335/net13	I0/I3335/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3332/T4	vss	I0/I3332/net13	I0/I3332/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3310/T4	vss	I0/I3310/net13	I0/I3310/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3323/T3	I0/I3323/net049	net946	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3313/T3	I0/I3313/net049	net945	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3339/T3	I0/I3339/net049	net944	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3333/T3	I0/I3333/net049	net943	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3319/T3	I0/I3319/net049	net942	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3312/T3	I0/I3312/net049	net941	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3335/T3	I0/I3335/net049	net940	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3332/T3	I0/I3332/net049	net939	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3310/T3	I0/I3310/net049	net938	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3355/T4	vss	I0/I3355/net13	I0/I3355/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3345/T4	vss	I0/I3345/net13	I0/I3345/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3355/T5	I0/I3355/net13	I0/I3355/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3345/T5	I0/I3345/net13	I0/I3345/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3355/T2	BL14	net946	I0/I3355/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3345/T2	BL14	net945	I0/I3345/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3371/T4	vss	I0/I3371/net13	I0/I3371/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3365/T4	vss	I0/I3365/net13	I0/I3365/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3371/T5	I0/I3371/net13	I0/I3371/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3365/T5	I0/I3365/net13	I0/I3365/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3371/T2	BL14	net944	I0/I3371/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3365/T2	BL14	net943	I0/I3365/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3351/T4	vss	I0/I3351/net13	I0/I3351/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3351/T5	I0/I3351/net13	I0/I3351/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3351/T2	BL14	net942	I0/I3351/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3344/T4	vss	I0/I3344/net13	I0/I3344/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3367/T4	vss	I0/I3367/net13	I0/I3367/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3344/T5	I0/I3344/net13	I0/I3344/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3367/T5	I0/I3367/net13	I0/I3367/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3344/T2	BL14	net941	I0/I3344/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3367/T2	BL14	net940	I0/I3367/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3364/T4	vss	I0/I3364/net13	I0/I3364/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3342/T4	vss	I0/I3342/net13	I0/I3342/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3364/T5	I0/I3364/net13	I0/I3364/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3342/T5	I0/I3342/net13	I0/I3342/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3364/T2	BL14	net939	I0/I3364/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3342/T2	BL14	net938	I0/I3342/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3355/T3	I0/I3355/net049	net946	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3345/T3	I0/I3345/net049	net945	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3371/T3	I0/I3371/net049	net944	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3365/T3	I0/I3365/net049	net943	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3351/T3	I0/I3351/net049	net942	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3344/T3	I0/I3344/net049	net941	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3367/T3	I0/I3367/net049	net940	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3364/T3	I0/I3364/net049	net939	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3342/T3	I0/I3342/net049	net938	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3387/T2	BL15	net946	I0/I3387/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3377/T2	BL15	net945	I0/I3377/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3403/T2	BL15	net944	I0/I3403/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3397/T2	BL15	net943	I0/I3397/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3383/T2	BL15	net942	I0/I3383/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3376/T2	BL15	net941	I0/I3376/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3399/T2	BL15	net940	I0/I3399/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3396/T2	BL15	net939	I0/I3396/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3374/T2	BL15	net938	I0/I3374/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3387/T5	I0/I3387/net13	I0/I3387/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3377/T5	I0/I3377/net13	I0/I3377/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3403/T5	I0/I3403/net13	I0/I3403/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3397/T5	I0/I3397/net13	I0/I3397/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3383/T5	I0/I3383/net13	I0/I3383/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3376/T5	I0/I3376/net13	I0/I3376/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3399/T5	I0/I3399/net13	I0/I3399/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3396/T5	I0/I3396/net13	I0/I3396/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3374/T5	I0/I3374/net13	I0/I3374/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3387/T4	vss	I0/I3387/net13	I0/I3387/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3377/T4	vss	I0/I3377/net13	I0/I3377/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3403/T4	vss	I0/I3403/net13	I0/I3403/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3397/T4	vss	I0/I3397/net13	I0/I3397/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3383/T4	vss	I0/I3383/net13	I0/I3383/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3376/T4	vss	I0/I3376/net13	I0/I3376/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3399/T4	vss	I0/I3399/net13	I0/I3399/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3396/T4	vss	I0/I3396/net13	I0/I3396/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3374/T4	vss	I0/I3374/net13	I0/I3374/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3387/T3	I0/I3387/net049	net946	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3377/T3	I0/I3377/net049	net945	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3403/T3	I0/I3403/net049	net944	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3397/T3	I0/I3397/net049	net943	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3383/T3	I0/I3383/net049	net942	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3376/T3	I0/I3376/net049	net941	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3399/T3	I0/I3399/net049	net940	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3396/T3	I0/I3396/net049	net939	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3374/T3	I0/I3374/net049	net938	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3099/T2	BL8	net946	I0/I3099/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3089/T2	BL8	net945	I0/I3089/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3115/T2	BL8	net944	I0/I3115/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3109/T2	BL8	net943	I0/I3109/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3095/T2	BL8	net942	I0/I3095/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3088/T2	BL8	net941	I0/I3088/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3111/T2	BL8	net940	I0/I3111/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3108/T2	BL8	net939	I0/I3108/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3086/T2	BL8	net938	I0/I3086/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3471/T3	I0/I3471/net049	net937	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3471/T4	vss	I0/I3471/net13	I0/I3471/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3471/T5	I0/I3471/net13	I0/I3471/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3471/T2	BL18	net937	I0/I3471/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3439/T3	I0/I3439/net049	net937	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3439/T4	vss	I0/I3439/net13	I0/I3439/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3439/T5	I0/I3439/net13	I0/I3439/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3279/T4	vss	I0/I3279/net13	I0/I3279/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3279/T5	I0/I3279/net13	I0/I3279/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3279/T2	BL12	net937	I0/I3279/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3503/T3	I0/I3503/net049	net937	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3503/T4	vss	I0/I3503/net13	I0/I3503/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3503/T5	I0/I3503/net13	I0/I3503/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3503/T2	BL19	net937	I0/I3503/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3279/T3	I0/I3279/net049	net937	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3343/T4	vss	I0/I3343/net13	I0/I3343/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3343/T5	I0/I3343/net13	I0/I3343/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3343/T2	BL14	net937	I0/I3343/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3311/T3	I0/I3311/net049	net937	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3311/T4	vss	I0/I3311/net13	I0/I3311/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3311/T5	I0/I3311/net13	I0/I3311/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3311/T2	BL13	net937	I0/I3311/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3087/T2	BL8	net937	I0/I3087/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3375/T3	I0/I3375/net049	net937	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3375/T4	vss	I0/I3375/net13	I0/I3375/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3375/T5	I0/I3375/net13	I0/I3375/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3375/T2	BL15	net937	I0/I3375/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3343/T3	I0/I3343/net049	net937	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3446/T3	I0/I3446/net049	net936	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3448/T3	I0/I3448/net049	net935	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3446/T4	vss	I0/I3446/net13	I0/I3446/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3448/T4	vss	I0/I3448/net13	I0/I3448/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3446/T5	I0/I3446/net13	I0/I3446/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3448/T5	I0/I3448/net13	I0/I3448/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3454/T3	I0/I3454/net049	net934	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3456/T3	I0/I3456/net049	net933	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3454/T4	vss	I0/I3454/net13	I0/I3454/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3456/T4	vss	I0/I3456/net13	I0/I3456/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3454/T5	I0/I3454/net13	I0/I3454/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3456/T5	I0/I3456/net13	I0/I3456/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3445/T3	I0/I3445/net049	net932	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3445/T4	vss	I0/I3445/net13	I0/I3445/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3445/T5	I0/I3445/net13	I0/I3445/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3459/T3	I0/I3459/net049	net931	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3453/T3	I0/I3453/net049	net930	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3459/T4	vss	I0/I3459/net13	I0/I3459/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3453/T4	vss	I0/I3453/net13	I0/I3453/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3459/T5	I0/I3459/net13	I0/I3459/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3453/T5	I0/I3453/net13	I0/I3453/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3457/T3	I0/I3457/net049	net929	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3469/T3	I0/I3469/net049	net928	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3457/T4	vss	I0/I3457/net13	I0/I3457/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3469/T4	vss	I0/I3469/net13	I0/I3469/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3457/T5	I0/I3457/net13	I0/I3457/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3469/T5	I0/I3469/net13	I0/I3469/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3478/T2	BL18	net936	I0/I3478/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3480/T2	BL18	net935	I0/I3480/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3486/T2	BL18	net934	I0/I3486/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3488/T2	BL18	net933	I0/I3488/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3477/T2	BL18	net932	I0/I3477/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3491/T2	BL18	net931	I0/I3491/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3485/T2	BL18	net930	I0/I3485/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3489/T2	BL18	net929	I0/I3489/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3501/T2	BL18	net928	I0/I3501/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3478/T5	I0/I3478/net13	I0/I3478/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3480/T5	I0/I3480/net13	I0/I3480/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3486/T5	I0/I3486/net13	I0/I3486/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3488/T5	I0/I3488/net13	I0/I3488/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3477/T5	I0/I3477/net13	I0/I3477/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3491/T5	I0/I3491/net13	I0/I3491/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3485/T5	I0/I3485/net13	I0/I3485/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3489/T5	I0/I3489/net13	I0/I3489/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3501/T5	I0/I3501/net13	I0/I3501/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3478/T4	vss	I0/I3478/net13	I0/I3478/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3480/T4	vss	I0/I3480/net13	I0/I3480/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3486/T4	vss	I0/I3486/net13	I0/I3486/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3488/T4	vss	I0/I3488/net13	I0/I3488/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3477/T4	vss	I0/I3477/net13	I0/I3477/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3491/T4	vss	I0/I3491/net13	I0/I3491/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3485/T4	vss	I0/I3485/net13	I0/I3485/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3489/T4	vss	I0/I3489/net13	I0/I3489/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3501/T4	vss	I0/I3501/net13	I0/I3501/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3478/T3	I0/I3478/net049	net936	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3480/T3	I0/I3480/net049	net935	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3486/T3	I0/I3486/net049	net934	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3488/T3	I0/I3488/net049	net933	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3477/T3	I0/I3477/net049	net932	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3491/T3	I0/I3491/net049	net931	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3485/T3	I0/I3485/net049	net930	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3489/T3	I0/I3489/net049	net929	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3501/T3	I0/I3501/net049	net928	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3510/T2	BL19	net936	I0/I3510/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3512/T2	BL19	net935	I0/I3512/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3518/T2	BL19	net934	I0/I3518/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3520/T2	BL19	net933	I0/I3520/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3509/T2	BL19	net932	I0/I3509/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3523/T2	BL19	net931	I0/I3523/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3517/T2	BL19	net930	I0/I3517/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3521/T2	BL19	net929	I0/I3521/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3533/T2	BL19	net928	I0/I3533/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3510/T5	I0/I3510/net13	I0/I3510/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3512/T5	I0/I3512/net13	I0/I3512/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3518/T5	I0/I3518/net13	I0/I3518/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3520/T5	I0/I3520/net13	I0/I3520/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3509/T5	I0/I3509/net13	I0/I3509/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3523/T5	I0/I3523/net13	I0/I3523/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3517/T5	I0/I3517/net13	I0/I3517/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3521/T5	I0/I3521/net13	I0/I3521/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3533/T5	I0/I3533/net13	I0/I3533/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3510/T4	vss	I0/I3510/net13	I0/I3510/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3512/T4	vss	I0/I3512/net13	I0/I3512/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3518/T4	vss	I0/I3518/net13	I0/I3518/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3520/T4	vss	I0/I3520/net13	I0/I3520/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3509/T4	vss	I0/I3509/net13	I0/I3509/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3523/T4	vss	I0/I3523/net13	I0/I3523/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3517/T4	vss	I0/I3517/net13	I0/I3517/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3521/T4	vss	I0/I3521/net13	I0/I3521/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3533/T4	vss	I0/I3533/net13	I0/I3533/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3510/T3	I0/I3510/net049	net936	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3512/T3	I0/I3512/net049	net935	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3518/T3	I0/I3518/net049	net934	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3520/T3	I0/I3520/net049	net933	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3509/T3	I0/I3509/net049	net932	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3523/T3	I0/I3523/net049	net931	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3517/T3	I0/I3517/net049	net930	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3521/T3	I0/I3521/net049	net929	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3533/T3	I0/I3533/net049	net928	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3286/T4	vss	I0/I3286/net13	I0/I3286/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3288/T4	vss	I0/I3288/net13	I0/I3288/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3286/T5	I0/I3286/net13	I0/I3286/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3288/T5	I0/I3288/net13	I0/I3288/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3286/T2	BL12	net936	I0/I3286/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3288/T2	BL12	net935	I0/I3288/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3294/T4	vss	I0/I3294/net13	I0/I3294/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3296/T4	vss	I0/I3296/net13	I0/I3296/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3294/T5	I0/I3294/net13	I0/I3294/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3296/T5	I0/I3296/net13	I0/I3296/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3294/T2	BL12	net934	I0/I3294/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3296/T2	BL12	net933	I0/I3296/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3285/T4	vss	I0/I3285/net13	I0/I3285/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3285/T5	I0/I3285/net13	I0/I3285/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3285/T2	BL12	net932	I0/I3285/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3299/T4	vss	I0/I3299/net13	I0/I3299/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3293/T4	vss	I0/I3293/net13	I0/I3293/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3299/T5	I0/I3299/net13	I0/I3299/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3293/T5	I0/I3293/net13	I0/I3293/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3299/T2	BL12	net931	I0/I3299/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3293/T2	BL12	net930	I0/I3293/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3297/T4	vss	I0/I3297/net13	I0/I3297/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3309/T4	vss	I0/I3309/net13	I0/I3309/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3297/T5	I0/I3297/net13	I0/I3297/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3309/T5	I0/I3309/net13	I0/I3309/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3297/T2	BL12	net929	I0/I3297/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3309/T2	BL12	net928	I0/I3309/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3286/T3	I0/I3286/net049	net936	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3288/T3	I0/I3288/net049	net935	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3294/T3	I0/I3294/net049	net934	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3296/T3	I0/I3296/net049	net933	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3285/T3	I0/I3285/net049	net932	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3299/T3	I0/I3299/net049	net931	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3293/T3	I0/I3293/net049	net930	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3297/T3	I0/I3297/net049	net929	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3309/T3	I0/I3309/net049	net928	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3318/T2	BL13	net936	I0/I3318/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3320/T2	BL13	net935	I0/I3320/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3326/T2	BL13	net934	I0/I3326/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3328/T2	BL13	net933	I0/I3328/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3317/T2	BL13	net932	I0/I3317/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3331/T2	BL13	net931	I0/I3331/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3325/T2	BL13	net930	I0/I3325/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3329/T2	BL13	net929	I0/I3329/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3341/T2	BL13	net928	I0/I3341/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3318/T5	I0/I3318/net13	I0/I3318/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3320/T5	I0/I3320/net13	I0/I3320/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3326/T5	I0/I3326/net13	I0/I3326/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3328/T5	I0/I3328/net13	I0/I3328/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3317/T5	I0/I3317/net13	I0/I3317/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3331/T5	I0/I3331/net13	I0/I3331/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3325/T5	I0/I3325/net13	I0/I3325/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3329/T5	I0/I3329/net13	I0/I3329/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3341/T5	I0/I3341/net13	I0/I3341/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3318/T4	vss	I0/I3318/net13	I0/I3318/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3320/T4	vss	I0/I3320/net13	I0/I3320/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3326/T4	vss	I0/I3326/net13	I0/I3326/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3328/T4	vss	I0/I3328/net13	I0/I3328/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3317/T4	vss	I0/I3317/net13	I0/I3317/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3331/T4	vss	I0/I3331/net13	I0/I3331/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3325/T4	vss	I0/I3325/net13	I0/I3325/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3329/T4	vss	I0/I3329/net13	I0/I3329/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3341/T4	vss	I0/I3341/net13	I0/I3341/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3318/T3	I0/I3318/net049	net936	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3320/T3	I0/I3320/net049	net935	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3326/T3	I0/I3326/net049	net934	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3328/T3	I0/I3328/net049	net933	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3317/T3	I0/I3317/net049	net932	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3331/T3	I0/I3331/net049	net931	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3325/T3	I0/I3325/net049	net930	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3329/T3	I0/I3329/net049	net929	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3341/T3	I0/I3341/net049	net928	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3350/T4	vss	I0/I3350/net13	I0/I3350/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3352/T4	vss	I0/I3352/net13	I0/I3352/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3350/T5	I0/I3350/net13	I0/I3350/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3352/T5	I0/I3352/net13	I0/I3352/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3350/T2	BL14	net936	I0/I3350/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3352/T2	BL14	net935	I0/I3352/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3358/T4	vss	I0/I3358/net13	I0/I3358/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3360/T4	vss	I0/I3360/net13	I0/I3360/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3358/T5	I0/I3358/net13	I0/I3358/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3360/T5	I0/I3360/net13	I0/I3360/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3358/T2	BL14	net934	I0/I3358/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3360/T2	BL14	net933	I0/I3360/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3349/T4	vss	I0/I3349/net13	I0/I3349/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3349/T5	I0/I3349/net13	I0/I3349/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3349/T2	BL14	net932	I0/I3349/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3363/T4	vss	I0/I3363/net13	I0/I3363/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3357/T4	vss	I0/I3357/net13	I0/I3357/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3363/T5	I0/I3363/net13	I0/I3363/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3357/T5	I0/I3357/net13	I0/I3357/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3363/T2	BL14	net931	I0/I3363/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3357/T2	BL14	net930	I0/I3357/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3361/T4	vss	I0/I3361/net13	I0/I3361/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3373/T4	vss	I0/I3373/net13	I0/I3373/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3361/T5	I0/I3361/net13	I0/I3361/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3373/T5	I0/I3373/net13	I0/I3373/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3361/T2	BL14	net929	I0/I3361/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3373/T2	BL14	net928	I0/I3373/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3350/T3	I0/I3350/net049	net936	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3352/T3	I0/I3352/net049	net935	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3358/T3	I0/I3358/net049	net934	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3360/T3	I0/I3360/net049	net933	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3349/T3	I0/I3349/net049	net932	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3363/T3	I0/I3363/net049	net931	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3357/T3	I0/I3357/net049	net930	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3361/T3	I0/I3361/net049	net929	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3373/T3	I0/I3373/net049	net928	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3382/T2	BL15	net936	I0/I3382/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3384/T2	BL15	net935	I0/I3384/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3390/T2	BL15	net934	I0/I3390/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3392/T2	BL15	net933	I0/I3392/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3381/T2	BL15	net932	I0/I3381/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3395/T2	BL15	net931	I0/I3395/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3389/T2	BL15	net930	I0/I3389/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3393/T2	BL15	net929	I0/I3393/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3405/T2	BL15	net928	I0/I3405/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3382/T5	I0/I3382/net13	I0/I3382/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3384/T5	I0/I3384/net13	I0/I3384/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3390/T5	I0/I3390/net13	I0/I3390/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3392/T5	I0/I3392/net13	I0/I3392/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3381/T5	I0/I3381/net13	I0/I3381/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3395/T5	I0/I3395/net13	I0/I3395/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3389/T5	I0/I3389/net13	I0/I3389/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3393/T5	I0/I3393/net13	I0/I3393/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3405/T5	I0/I3405/net13	I0/I3405/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3382/T4	vss	I0/I3382/net13	I0/I3382/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3384/T4	vss	I0/I3384/net13	I0/I3384/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3390/T4	vss	I0/I3390/net13	I0/I3390/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3392/T4	vss	I0/I3392/net13	I0/I3392/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3381/T4	vss	I0/I3381/net13	I0/I3381/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3395/T4	vss	I0/I3395/net13	I0/I3395/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3389/T4	vss	I0/I3389/net13	I0/I3389/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3393/T4	vss	I0/I3393/net13	I0/I3393/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3405/T4	vss	I0/I3405/net13	I0/I3405/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3382/T3	I0/I3382/net049	net936	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3384/T3	I0/I3384/net049	net935	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3390/T3	I0/I3390/net049	net934	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3392/T3	I0/I3392/net049	net933	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3381/T3	I0/I3381/net049	net932	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3395/T3	I0/I3395/net049	net931	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3389/T3	I0/I3389/net049	net930	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3393/T3	I0/I3393/net049	net929	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3405/T3	I0/I3405/net049	net928	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3094/T2	BL8	net936	I0/I3094/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3096/T2	BL8	net935	I0/I3096/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3102/T2	BL8	net934	I0/I3102/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3104/T2	BL8	net933	I0/I3104/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3093/T2	BL8	net932	I0/I3093/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3107/T2	BL8	net931	I0/I3107/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3101/T2	BL8	net930	I0/I3101/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3105/T2	BL8	net929	I0/I3105/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3117/T2	BL8	net928	I0/I3117/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3487/T3	I0/I3487/net049	net927	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3487/T4	vss	I0/I3487/net13	I0/I3487/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3487/T5	I0/I3487/net13	I0/I3487/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3487/T2	BL18	net927	I0/I3487/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3455/T3	I0/I3455/net049	net927	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3455/T4	vss	I0/I3455/net13	I0/I3455/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3455/T5	I0/I3455/net13	I0/I3455/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3295/T4	vss	I0/I3295/net13	I0/I3295/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3295/T5	I0/I3295/net13	I0/I3295/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3295/T2	BL12	net927	I0/I3295/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3519/T3	I0/I3519/net049	net927	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3519/T4	vss	I0/I3519/net13	I0/I3519/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3519/T5	I0/I3519/net13	I0/I3519/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3519/T2	BL19	net927	I0/I3519/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3295/T3	I0/I3295/net049	net927	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3359/T4	vss	I0/I3359/net13	I0/I3359/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3359/T5	I0/I3359/net13	I0/I3359/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3359/T2	BL14	net927	I0/I3359/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3327/T3	I0/I3327/net049	net927	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3327/T4	vss	I0/I3327/net13	I0/I3327/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3327/T5	I0/I3327/net13	I0/I3327/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3327/T2	BL13	net927	I0/I3327/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3103/T2	BL8	net927	I0/I3103/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3391/T3	I0/I3391/net049	net927	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3391/T4	vss	I0/I3391/net13	I0/I3391/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3391/T5	I0/I3391/net13	I0/I3391/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3391/T2	BL15	net927	I0/I3391/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3359/T3	I0/I3359/net049	net927	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3498/T3	I0/I3498/net049	net926	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3498/T4	vss	I0/I3498/net13	I0/I3498/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3498/T5	I0/I3498/net13	I0/I3498/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3498/T2	BL18	net926	I0/I3498/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3466/T3	I0/I3466/net049	net926	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3466/T4	vss	I0/I3466/net13	I0/I3466/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3466/T5	I0/I3466/net13	I0/I3466/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3306/T4	vss	I0/I3306/net13	I0/I3306/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3306/T5	I0/I3306/net13	I0/I3306/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3306/T2	BL12	net926	I0/I3306/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3530/T3	I0/I3530/net049	net926	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3530/T4	vss	I0/I3530/net13	I0/I3530/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3530/T5	I0/I3530/net13	I0/I3530/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3530/T2	BL19	net926	I0/I3530/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3306/T3	I0/I3306/net049	net926	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3370/T4	vss	I0/I3370/net13	I0/I3370/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3370/T5	I0/I3370/net13	I0/I3370/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3370/T2	BL14	net926	I0/I3370/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3338/T3	I0/I3338/net049	net926	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3338/T4	vss	I0/I3338/net13	I0/I3338/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3338/T5	I0/I3338/net13	I0/I3338/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3338/T2	BL13	net926	I0/I3338/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3114/T2	BL8	net926	I0/I3114/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3402/T3	I0/I3402/net049	net926	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3402/T4	vss	I0/I3402/net13	I0/I3402/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3402/T5	I0/I3402/net13	I0/I3402/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3402/T2	BL15	net926	I0/I3402/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3370/T3	I0/I3370/net049	net926	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3497/T3	I0/I3497/net049	net925	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3497/T4	vss	I0/I3497/net13	I0/I3497/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3497/T5	I0/I3497/net13	I0/I3497/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3497/T2	BL18	net925	I0/I3497/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3465/T3	I0/I3465/net049	net925	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3465/T4	vss	I0/I3465/net13	I0/I3465/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3465/T5	I0/I3465/net13	I0/I3465/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3305/T4	vss	I0/I3305/net13	I0/I3305/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3305/T5	I0/I3305/net13	I0/I3305/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3305/T2	BL12	net925	I0/I3305/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3529/T3	I0/I3529/net049	net925	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3529/T4	vss	I0/I3529/net13	I0/I3529/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3529/T5	I0/I3529/net13	I0/I3529/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3529/T2	BL19	net925	I0/I3529/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3305/T3	I0/I3305/net049	net925	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3369/T4	vss	I0/I3369/net13	I0/I3369/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3369/T5	I0/I3369/net13	I0/I3369/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3369/T2	BL14	net925	I0/I3369/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3337/T3	I0/I3337/net049	net925	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3337/T4	vss	I0/I3337/net13	I0/I3337/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3337/T5	I0/I3337/net13	I0/I3337/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3337/T2	BL13	net925	I0/I3337/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3113/T2	BL8	net925	I0/I3113/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3401/T3	I0/I3401/net049	net925	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3401/T4	vss	I0/I3401/net13	I0/I3401/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3401/T5	I0/I3401/net13	I0/I3401/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3401/T2	BL15	net925	I0/I3401/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3369/T3	I0/I3369/net049	net925	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3474/T3	I0/I3474/net049	net924	BL18bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3474/T4	vss	I0/I3474/net13	I0/I3474/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3474/T5	I0/I3474/net13	I0/I3474/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3474/T2	BL18	net924	I0/I3474/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3442/T3	I0/I3442/net049	net924	BL17bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3442/T4	vss	I0/I3442/net13	I0/I3442/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3442/T5	I0/I3442/net13	I0/I3442/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3282/T4	vss	I0/I3282/net13	I0/I3282/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3282/T5	I0/I3282/net13	I0/I3282/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3282/T2	BL12	net924	I0/I3282/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3506/T3	I0/I3506/net049	net924	BL19bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3506/T4	vss	I0/I3506/net13	I0/I3506/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3506/T5	I0/I3506/net13	I0/I3506/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3506/T2	BL19	net924	I0/I3506/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3282/T3	I0/I3282/net049	net924	BL12bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3346/T4	vss	I0/I3346/net13	I0/I3346/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3346/T5	I0/I3346/net13	I0/I3346/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3346/T2	BL14	net924	I0/I3346/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3314/T3	I0/I3314/net049	net924	BL13bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3314/T4	vss	I0/I3314/net13	I0/I3314/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3314/T5	I0/I3314/net13	I0/I3314/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3314/T2	BL13	net924	I0/I3314/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3090/T2	BL8	net924	I0/I3090/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3378/T3	I0/I3378/net049	net924	BL15bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3378/T4	vss	I0/I3378/net13	I0/I3378/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3378/T5	I0/I3378/net13	I0/I3378/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3378/T2	BL15	net924	I0/I3378/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3346/T3	I0/I3346/net049	net924	BL14bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI66/T1	p4bar	y1	BL12bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI67/T1	BL12	y1	p4	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI68/T1	p5bar	y4	BL19bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI69/T1	BL19	y4	p5	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI70/T1	p5bar	y3	BL18bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI71/T1	BL18	y3	p5	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI72/T1	p5bar	y2	BL17bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI59/T1	BL8	y1	net740	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI60/T1	p4bar	y4	BL15bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI61/T1	BL15	y4	p4	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI62/T1	p4bar	y3	BL14bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI63/T1	BL14	y3	p4	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI64/T1	p4bar	y2	BL13bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI65/T1	BL13	y2	p4	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T3	I3/net20	net741	I3/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T4	vss	vdd	I3/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T8	vss	I3/net20	I3/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T7	data2	I3/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T11	I25/net23	data2	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T16	I25/net15	net680	net740	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T17	vss	I25/net23	I25/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T19	I25/net7	net740	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T18	net741	net680	I25/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T8	vss	I2/net20	I2/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T7	data1	I2/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T11	I24/net23	data1	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T16	I24/net15	net680	net262	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T17	vss	I24/net23	I24/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T19	I24/net7	net262	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T18	net256	net680	I24/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T2	I3/net23	net740	I3/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T20	I30/net17	I30/net49	vss	vss	nfet	L=0.12U
+ W=0.64U
+ AD=0.2048P	AS=0.2048P	PD=1.92U	PS=1.92U
+ wt=6.4e-07 wf=6.4e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.68e-14 panw7=1.008e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.369748 nrd=0.369748 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI30/T3	I30/net49	wr	vss	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=4.32e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI30/T0	I30/net61	wr	vss	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=4.32e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI30/T14	I30/net57	I30/net61	vss	vss	nfet	L=0.12U
+ W=1.22U
+ AD=0.3904P	AS=0.3904P	PD=3.08U	PS=3.08U
+ wt=1.22e-06 wf=1.22e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.04e-14 panw7=1.464e-13 panw10=1.14e-13 nrs=0.187234 nrd=0.187234 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI30/T19	net681	I30/net57	vss	vss	nfet	L=0.12U
+ W=4.5U
+ AD=1.44P	AS=1.44P	PD=9.64U	PS=9.64U
+ wt=4.5e-06 wf=4.5e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=4.368e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0493827 nrd=0.0493827 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3100/T3	I0/I3100/net049	net955	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3092/T3	I0/I3092/net049	net954	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3100/T4	vss	I0/I3100/net13	I0/I3100/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3092/T4	vss	I0/I3092/net13	I0/I3092/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3100/T5	I0/I3100/net13	I0/I3100/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3092/T5	I0/I3092/net13	I0/I3092/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3091/T3	I0/I3091/net049	net953	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3116/T3	I0/I3116/net049	net952	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3091/T4	vss	I0/I3091/net13	I0/I3091/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3116/T4	vss	I0/I3116/net13	I0/I3116/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3091/T5	I0/I3091/net13	I0/I3091/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3116/T5	I0/I3116/net13	I0/I3116/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3097/T3	I0/I3097/net049	net951	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3097/T4	vss	I0/I3097/net13	I0/I3097/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3097/T5	I0/I3097/net13	I0/I3097/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3112/T3	I0/I3112/net049	net950	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3110/T3	I0/I3110/net049	net949	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3112/T4	vss	I0/I3112/net13	I0/I3112/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3110/T4	vss	I0/I3110/net13	I0/I3110/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3112/T5	I0/I3112/net13	I0/I3112/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3110/T5	I0/I3110/net13	I0/I3110/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3106/T3	I0/I3106/net049	net948	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3098/T3	I0/I3098/net049	net947	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3106/T4	vss	I0/I3106/net13	I0/I3106/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3098/T4	vss	I0/I3098/net13	I0/I3098/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3106/T5	I0/I3106/net13	I0/I3106/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3098/T5	I0/I3098/net13	I0/I3098/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3132/T2	BL9	net955	I0/I3132/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3124/T2	BL9	net954	I0/I3124/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3123/T2	BL9	net953	I0/I3123/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3148/T2	BL9	net952	I0/I3148/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3129/T2	BL9	net951	I0/I3129/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3144/T2	BL9	net950	I0/I3144/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3142/T2	BL9	net949	I0/I3142/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3138/T2	BL9	net948	I0/I3138/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3130/T2	BL9	net947	I0/I3130/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3132/T5	I0/I3132/net13	I0/I3132/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3124/T5	I0/I3124/net13	I0/I3124/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3123/T5	I0/I3123/net13	I0/I3123/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3148/T5	I0/I3148/net13	I0/I3148/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3129/T5	I0/I3129/net13	I0/I3129/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3144/T5	I0/I3144/net13	I0/I3144/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3142/T5	I0/I3142/net13	I0/I3142/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3138/T5	I0/I3138/net13	I0/I3138/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3130/T5	I0/I3130/net13	I0/I3130/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3132/T4	vss	I0/I3132/net13	I0/I3132/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3124/T4	vss	I0/I3124/net13	I0/I3124/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3123/T4	vss	I0/I3123/net13	I0/I3123/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3148/T4	vss	I0/I3148/net13	I0/I3148/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3129/T4	vss	I0/I3129/net13	I0/I3129/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3144/T4	vss	I0/I3144/net13	I0/I3144/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3142/T4	vss	I0/I3142/net13	I0/I3142/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3138/T4	vss	I0/I3138/net13	I0/I3138/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3130/T4	vss	I0/I3130/net13	I0/I3130/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3132/T3	I0/I3132/net049	net955	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3124/T3	I0/I3124/net049	net954	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3123/T3	I0/I3123/net049	net953	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3148/T3	I0/I3148/net049	net952	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3129/T3	I0/I3129/net049	net951	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3144/T3	I0/I3144/net049	net950	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3142/T3	I0/I3142/net049	net949	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3138/T3	I0/I3138/net049	net948	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3130/T3	I0/I3130/net049	net947	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3164/T2	BL10	net955	I0/I3164/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3156/T2	BL10	net954	I0/I3156/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3155/T2	BL10	net953	I0/I3155/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3180/T2	BL10	net952	I0/I3180/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3161/T2	BL10	net951	I0/I3161/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3176/T2	BL10	net950	I0/I3176/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3174/T2	BL10	net949	I0/I3174/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3170/T2	BL10	net948	I0/I3170/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3162/T2	BL10	net947	I0/I3162/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3164/T5	I0/I3164/net13	I0/I3164/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3156/T5	I0/I3156/net13	I0/I3156/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3155/T5	I0/I3155/net13	I0/I3155/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3180/T5	I0/I3180/net13	I0/I3180/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3161/T5	I0/I3161/net13	I0/I3161/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3176/T5	I0/I3176/net13	I0/I3176/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3174/T5	I0/I3174/net13	I0/I3174/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3170/T5	I0/I3170/net13	I0/I3170/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3162/T5	I0/I3162/net13	I0/I3162/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3164/T4	vss	I0/I3164/net13	I0/I3164/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3156/T4	vss	I0/I3156/net13	I0/I3156/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3155/T4	vss	I0/I3155/net13	I0/I3155/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3180/T4	vss	I0/I3180/net13	I0/I3180/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3161/T4	vss	I0/I3161/net13	I0/I3161/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3176/T4	vss	I0/I3176/net13	I0/I3176/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3174/T4	vss	I0/I3174/net13	I0/I3174/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3170/T4	vss	I0/I3170/net13	I0/I3170/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3162/T4	vss	I0/I3162/net13	I0/I3162/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3164/T3	I0/I3164/net049	net955	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3156/T3	I0/I3156/net049	net954	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3155/T3	I0/I3155/net049	net953	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3180/T3	I0/I3180/net049	net952	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3161/T3	I0/I3161/net049	net951	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3176/T3	I0/I3176/net049	net950	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3174/T3	I0/I3174/net049	net949	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3170/T3	I0/I3170/net049	net948	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3162/T3	I0/I3162/net049	net947	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3196/T4	vss	I0/I3196/net13	I0/I3196/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3188/T4	vss	I0/I3188/net13	I0/I3188/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3196/T5	I0/I3196/net13	I0/I3196/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3188/T5	I0/I3188/net13	I0/I3188/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3196/T2	BL11	net955	I0/I3196/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3188/T2	BL11	net954	I0/I3188/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3187/T4	vss	I0/I3187/net13	I0/I3187/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3212/T4	vss	I0/I3212/net13	I0/I3212/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3187/T5	I0/I3187/net13	I0/I3187/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3212/T5	I0/I3212/net13	I0/I3212/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3187/T2	BL11	net953	I0/I3187/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3212/T2	BL11	net952	I0/I3212/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3193/T4	vss	I0/I3193/net13	I0/I3193/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3193/T5	I0/I3193/net13	I0/I3193/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3193/T2	BL11	net951	I0/I3193/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3208/T4	vss	I0/I3208/net13	I0/I3208/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3206/T4	vss	I0/I3206/net13	I0/I3206/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3208/T5	I0/I3208/net13	I0/I3208/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3206/T5	I0/I3206/net13	I0/I3206/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3208/T2	BL11	net950	I0/I3208/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3206/T2	BL11	net949	I0/I3206/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3202/T4	vss	I0/I3202/net13	I0/I3202/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3194/T4	vss	I0/I3194/net13	I0/I3194/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3202/T5	I0/I3202/net13	I0/I3202/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3194/T5	I0/I3194/net13	I0/I3194/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3202/T2	BL11	net948	I0/I3202/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3194/T2	BL11	net947	I0/I3194/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3196/T3	I0/I3196/net049	net955	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3188/T3	I0/I3188/net049	net954	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3187/T3	I0/I3187/net049	net953	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3212/T3	I0/I3212/net049	net952	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3193/T3	I0/I3193/net049	net951	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3208/T3	I0/I3208/net049	net950	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3206/T3	I0/I3206/net049	net949	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3202/T3	I0/I3202/net049	net948	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3194/T3	I0/I3194/net049	net947	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I107/T2	BL4	net955	I0/I107/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I115/T2	BL4	net954	I0/I115/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I116/T2	BL4	net953	I0/I116/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I91/T2	BL4	net952	I0/I91/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I110/T2	BL4	net951	I0/I110/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I95/T2	BL4	net950	I0/I95/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I97/T2	BL4	net949	I0/I97/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I101/T2	BL4	net948	I0/I101/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I109/T2	BL4	net947	I0/I109/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I107/T5	I0/I107/net13	I0/I107/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I115/T5	I0/I115/net13	I0/I115/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I116/T5	I0/I116/net13	I0/I116/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I91/T5	I0/I91/net13	I0/I91/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I110/T5	I0/I110/net13	I0/I110/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I95/T5	I0/I95/net13	I0/I95/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I97/T5	I0/I97/net13	I0/I97/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I101/T5	I0/I101/net13	I0/I101/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I109/T5	I0/I109/net13	I0/I109/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I107/T4	vss	I0/I107/net13	I0/I107/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I115/T4	vss	I0/I115/net13	I0/I115/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I116/T4	vss	I0/I116/net13	I0/I116/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I91/T4	vss	I0/I91/net13	I0/I91/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I110/T4	vss	I0/I110/net13	I0/I110/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I95/T4	vss	I0/I95/net13	I0/I95/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I97/T4	vss	I0/I97/net13	I0/I97/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I101/T4	vss	I0/I101/net13	I0/I101/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I109/T4	vss	I0/I109/net13	I0/I109/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I107/T3	I0/I107/net049	net955	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I115/T3	I0/I115/net049	net954	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I116/T3	I0/I116/net049	net953	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I91/T3	I0/I91/net049	net952	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I110/T3	I0/I110/net049	net951	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I95/T3	I0/I95/net049	net950	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I97/T3	I0/I97/net049	net949	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I101/T3	I0/I101/net049	net948	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I109/T3	I0/I109/net049	net947	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3004/T4	vss	I0/I3004/net13	I0/I3004/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2996/T4	vss	I0/I2996/net13	I0/I2996/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3004/T5	I0/I3004/net13	I0/I3004/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2996/T5	I0/I2996/net13	I0/I2996/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3004/T2	BL5	net955	I0/I3004/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2996/T2	BL5	net954	I0/I2996/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2995/T4	vss	I0/I2995/net13	I0/I2995/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3020/T4	vss	I0/I3020/net13	I0/I3020/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2995/T5	I0/I2995/net13	I0/I2995/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3020/T5	I0/I3020/net13	I0/I3020/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2995/T2	BL5	net953	I0/I2995/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3020/T2	BL5	net952	I0/I3020/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3001/T4	vss	I0/I3001/net13	I0/I3001/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3001/T5	I0/I3001/net13	I0/I3001/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3001/T2	BL5	net951	I0/I3001/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3016/T4	vss	I0/I3016/net13	I0/I3016/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3014/T4	vss	I0/I3014/net13	I0/I3014/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3016/T5	I0/I3016/net13	I0/I3016/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3014/T5	I0/I3014/net13	I0/I3014/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3016/T2	BL5	net950	I0/I3016/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3014/T2	BL5	net949	I0/I3014/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3010/T4	vss	I0/I3010/net13	I0/I3010/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3002/T4	vss	I0/I3002/net13	I0/I3002/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3010/T5	I0/I3010/net13	I0/I3010/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3002/T5	I0/I3002/net13	I0/I3002/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3010/T2	BL5	net948	I0/I3010/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3002/T2	BL5	net947	I0/I3002/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3004/T3	I0/I3004/net049	net955	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2996/T3	I0/I2996/net049	net954	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2995/T3	I0/I2995/net049	net953	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3020/T3	I0/I3020/net049	net952	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3001/T3	I0/I3001/net049	net951	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3016/T3	I0/I3016/net049	net950	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3014/T3	I0/I3014/net049	net949	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3010/T3	I0/I3010/net049	net948	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3002/T3	I0/I3002/net049	net947	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3036/T2	BL6	net955	I0/I3036/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3028/T2	BL6	net954	I0/I3028/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3027/T2	BL6	net953	I0/I3027/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3052/T2	BL6	net952	I0/I3052/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3033/T2	BL6	net951	I0/I3033/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3048/T2	BL6	net950	I0/I3048/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3046/T2	BL6	net949	I0/I3046/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3042/T2	BL6	net948	I0/I3042/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3034/T2	BL6	net947	I0/I3034/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3036/T5	I0/I3036/net13	I0/I3036/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3028/T5	I0/I3028/net13	I0/I3028/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3027/T5	I0/I3027/net13	I0/I3027/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3052/T5	I0/I3052/net13	I0/I3052/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3033/T5	I0/I3033/net13	I0/I3033/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3048/T5	I0/I3048/net13	I0/I3048/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3046/T5	I0/I3046/net13	I0/I3046/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3042/T5	I0/I3042/net13	I0/I3042/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3034/T5	I0/I3034/net13	I0/I3034/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3036/T4	vss	I0/I3036/net13	I0/I3036/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3028/T4	vss	I0/I3028/net13	I0/I3028/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3027/T4	vss	I0/I3027/net13	I0/I3027/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3052/T4	vss	I0/I3052/net13	I0/I3052/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3033/T4	vss	I0/I3033/net13	I0/I3033/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3048/T4	vss	I0/I3048/net13	I0/I3048/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3046/T4	vss	I0/I3046/net13	I0/I3046/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3042/T4	vss	I0/I3042/net13	I0/I3042/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3034/T4	vss	I0/I3034/net13	I0/I3034/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3036/T3	I0/I3036/net049	net955	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3028/T3	I0/I3028/net049	net954	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3027/T3	I0/I3027/net049	net953	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3052/T3	I0/I3052/net049	net952	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3033/T3	I0/I3033/net049	net951	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3048/T3	I0/I3048/net049	net950	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3046/T3	I0/I3046/net049	net949	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3042/T3	I0/I3042/net049	net948	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3034/T3	I0/I3034/net049	net947	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3068/T2	BL7	net955	I0/I3068/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3060/T2	BL7	net954	I0/I3060/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3059/T2	BL7	net953	I0/I3059/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3084/T2	BL7	net952	I0/I3084/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3065/T2	BL7	net951	I0/I3065/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3080/T2	BL7	net950	I0/I3080/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3078/T2	BL7	net949	I0/I3078/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3074/T2	BL7	net948	I0/I3074/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3066/T2	BL7	net947	I0/I3066/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3099/T3	I0/I3099/net049	net946	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3089/T3	I0/I3089/net049	net945	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3099/T4	vss	I0/I3099/net13	I0/I3099/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3089/T4	vss	I0/I3089/net13	I0/I3089/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3099/T5	I0/I3099/net13	I0/I3099/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3089/T5	I0/I3089/net13	I0/I3089/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3115/T3	I0/I3115/net049	net944	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3109/T3	I0/I3109/net049	net943	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3115/T4	vss	I0/I3115/net13	I0/I3115/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3109/T4	vss	I0/I3109/net13	I0/I3109/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3115/T5	I0/I3115/net13	I0/I3115/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3109/T5	I0/I3109/net13	I0/I3109/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3095/T3	I0/I3095/net049	net942	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3095/T4	vss	I0/I3095/net13	I0/I3095/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3095/T5	I0/I3095/net13	I0/I3095/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3088/T3	I0/I3088/net049	net941	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3111/T3	I0/I3111/net049	net940	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3088/T4	vss	I0/I3088/net13	I0/I3088/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3111/T4	vss	I0/I3111/net13	I0/I3111/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3088/T5	I0/I3088/net13	I0/I3088/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3111/T5	I0/I3111/net13	I0/I3111/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3108/T3	I0/I3108/net049	net939	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3086/T3	I0/I3086/net049	net938	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3108/T4	vss	I0/I3108/net13	I0/I3108/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3086/T4	vss	I0/I3086/net13	I0/I3086/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3108/T5	I0/I3108/net13	I0/I3108/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3086/T5	I0/I3086/net13	I0/I3086/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3131/T2	BL9	net946	I0/I3131/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3121/T2	BL9	net945	I0/I3121/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3147/T2	BL9	net944	I0/I3147/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3141/T2	BL9	net943	I0/I3141/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3127/T2	BL9	net942	I0/I3127/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3120/T2	BL9	net941	I0/I3120/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3143/T2	BL9	net940	I0/I3143/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3140/T2	BL9	net939	I0/I3140/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3118/T2	BL9	net938	I0/I3118/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3131/T5	I0/I3131/net13	I0/I3131/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3121/T5	I0/I3121/net13	I0/I3121/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3147/T5	I0/I3147/net13	I0/I3147/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3141/T5	I0/I3141/net13	I0/I3141/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3127/T5	I0/I3127/net13	I0/I3127/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3120/T5	I0/I3120/net13	I0/I3120/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3143/T5	I0/I3143/net13	I0/I3143/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3140/T5	I0/I3140/net13	I0/I3140/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3118/T5	I0/I3118/net13	I0/I3118/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3131/T4	vss	I0/I3131/net13	I0/I3131/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3121/T4	vss	I0/I3121/net13	I0/I3121/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3147/T4	vss	I0/I3147/net13	I0/I3147/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3141/T4	vss	I0/I3141/net13	I0/I3141/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3127/T4	vss	I0/I3127/net13	I0/I3127/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3120/T4	vss	I0/I3120/net13	I0/I3120/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3143/T4	vss	I0/I3143/net13	I0/I3143/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3140/T4	vss	I0/I3140/net13	I0/I3140/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3118/T4	vss	I0/I3118/net13	I0/I3118/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3131/T3	I0/I3131/net049	net946	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3121/T3	I0/I3121/net049	net945	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3147/T3	I0/I3147/net049	net944	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3141/T3	I0/I3141/net049	net943	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3127/T3	I0/I3127/net049	net942	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3120/T3	I0/I3120/net049	net941	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3143/T3	I0/I3143/net049	net940	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3140/T3	I0/I3140/net049	net939	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3118/T3	I0/I3118/net049	net938	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3163/T2	BL10	net946	I0/I3163/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3153/T2	BL10	net945	I0/I3153/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3179/T2	BL10	net944	I0/I3179/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3173/T2	BL10	net943	I0/I3173/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3159/T2	BL10	net942	I0/I3159/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3152/T2	BL10	net941	I0/I3152/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3175/T2	BL10	net940	I0/I3175/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3172/T2	BL10	net939	I0/I3172/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3150/T2	BL10	net938	I0/I3150/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3163/T5	I0/I3163/net13	I0/I3163/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3153/T5	I0/I3153/net13	I0/I3153/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3179/T5	I0/I3179/net13	I0/I3179/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3173/T5	I0/I3173/net13	I0/I3173/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3159/T5	I0/I3159/net13	I0/I3159/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3152/T5	I0/I3152/net13	I0/I3152/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3175/T5	I0/I3175/net13	I0/I3175/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3172/T5	I0/I3172/net13	I0/I3172/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3150/T5	I0/I3150/net13	I0/I3150/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3163/T4	vss	I0/I3163/net13	I0/I3163/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3153/T4	vss	I0/I3153/net13	I0/I3153/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3179/T4	vss	I0/I3179/net13	I0/I3179/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3173/T4	vss	I0/I3173/net13	I0/I3173/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3159/T4	vss	I0/I3159/net13	I0/I3159/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3152/T4	vss	I0/I3152/net13	I0/I3152/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3175/T4	vss	I0/I3175/net13	I0/I3175/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3172/T4	vss	I0/I3172/net13	I0/I3172/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3150/T4	vss	I0/I3150/net13	I0/I3150/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3163/T3	I0/I3163/net049	net946	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3153/T3	I0/I3153/net049	net945	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3179/T3	I0/I3179/net049	net944	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3173/T3	I0/I3173/net049	net943	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3159/T3	I0/I3159/net049	net942	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3152/T3	I0/I3152/net049	net941	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3175/T3	I0/I3175/net049	net940	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3172/T3	I0/I3172/net049	net939	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3150/T3	I0/I3150/net049	net938	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3195/T4	vss	I0/I3195/net13	I0/I3195/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3185/T4	vss	I0/I3185/net13	I0/I3185/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3195/T5	I0/I3195/net13	I0/I3195/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3185/T5	I0/I3185/net13	I0/I3185/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3195/T2	BL11	net946	I0/I3195/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3185/T2	BL11	net945	I0/I3185/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3211/T4	vss	I0/I3211/net13	I0/I3211/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3205/T4	vss	I0/I3205/net13	I0/I3205/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3211/T5	I0/I3211/net13	I0/I3211/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3205/T5	I0/I3205/net13	I0/I3205/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3211/T2	BL11	net944	I0/I3211/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3205/T2	BL11	net943	I0/I3205/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3191/T4	vss	I0/I3191/net13	I0/I3191/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3191/T5	I0/I3191/net13	I0/I3191/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3191/T2	BL11	net942	I0/I3191/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3184/T4	vss	I0/I3184/net13	I0/I3184/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3207/T4	vss	I0/I3207/net13	I0/I3207/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3184/T5	I0/I3184/net13	I0/I3184/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3207/T5	I0/I3207/net13	I0/I3207/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3184/T2	BL11	net941	I0/I3184/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3207/T2	BL11	net940	I0/I3207/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3204/T4	vss	I0/I3204/net13	I0/I3204/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3182/T4	vss	I0/I3182/net13	I0/I3182/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3204/T5	I0/I3204/net13	I0/I3204/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3182/T5	I0/I3182/net13	I0/I3182/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3204/T2	BL11	net939	I0/I3204/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3182/T2	BL11	net938	I0/I3182/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3195/T3	I0/I3195/net049	net946	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3185/T3	I0/I3185/net049	net945	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3211/T3	I0/I3211/net049	net944	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3205/T3	I0/I3205/net049	net943	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3191/T3	I0/I3191/net049	net942	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3184/T3	I0/I3184/net049	net941	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3207/T3	I0/I3207/net049	net940	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3204/T3	I0/I3204/net049	net939	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3182/T3	I0/I3182/net049	net938	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I108/T2	BL4	net946	I0/I108/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I118/T2	BL4	net945	I0/I118/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I92/T2	BL4	net944	I0/I92/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I98/T2	BL4	net943	I0/I98/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I112/T2	BL4	net942	I0/I112/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I119/T2	BL4	net941	I0/I119/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I96/T2	BL4	net940	I0/I96/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I99/T2	BL4	net939	I0/I99/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I121/T2	BL4	net938	I0/I121/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I108/T5	I0/I108/net13	I0/I108/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I118/T5	I0/I118/net13	I0/I118/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I92/T5	I0/I92/net13	I0/I92/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I98/T5	I0/I98/net13	I0/I98/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I112/T5	I0/I112/net13	I0/I112/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I119/T5	I0/I119/net13	I0/I119/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I96/T5	I0/I96/net13	I0/I96/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I99/T5	I0/I99/net13	I0/I99/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I121/T5	I0/I121/net13	I0/I121/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I108/T4	vss	I0/I108/net13	I0/I108/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I118/T4	vss	I0/I118/net13	I0/I118/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I92/T4	vss	I0/I92/net13	I0/I92/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I98/T4	vss	I0/I98/net13	I0/I98/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I112/T4	vss	I0/I112/net13	I0/I112/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I119/T4	vss	I0/I119/net13	I0/I119/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I96/T4	vss	I0/I96/net13	I0/I96/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I99/T4	vss	I0/I99/net13	I0/I99/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I121/T4	vss	I0/I121/net13	I0/I121/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I108/T3	I0/I108/net049	net946	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I118/T3	I0/I118/net049	net945	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I92/T3	I0/I92/net049	net944	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I98/T3	I0/I98/net049	net943	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I112/T3	I0/I112/net049	net942	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I119/T3	I0/I119/net049	net941	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I96/T3	I0/I96/net049	net940	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I99/T3	I0/I99/net049	net939	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I121/T3	I0/I121/net049	net938	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3003/T4	vss	I0/I3003/net13	I0/I3003/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2993/T4	vss	I0/I2993/net13	I0/I2993/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3003/T5	I0/I3003/net13	I0/I3003/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2993/T5	I0/I2993/net13	I0/I2993/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3003/T2	BL5	net946	I0/I3003/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2993/T2	BL5	net945	I0/I2993/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3019/T4	vss	I0/I3019/net13	I0/I3019/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3013/T4	vss	I0/I3013/net13	I0/I3013/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3019/T5	I0/I3019/net13	I0/I3019/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3013/T5	I0/I3013/net13	I0/I3013/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3019/T2	BL5	net944	I0/I3019/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3013/T2	BL5	net943	I0/I3013/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2999/T4	vss	I0/I2999/net13	I0/I2999/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2999/T5	I0/I2999/net13	I0/I2999/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2999/T2	BL5	net942	I0/I2999/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2992/T4	vss	I0/I2992/net13	I0/I2992/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3015/T4	vss	I0/I3015/net13	I0/I3015/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2992/T5	I0/I2992/net13	I0/I2992/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3015/T5	I0/I3015/net13	I0/I3015/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2992/T2	BL5	net941	I0/I2992/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3015/T2	BL5	net940	I0/I3015/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3012/T4	vss	I0/I3012/net13	I0/I3012/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2990/T4	vss	I0/I2990/net13	I0/I2990/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3012/T5	I0/I3012/net13	I0/I3012/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2990/T5	I0/I2990/net13	I0/I2990/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3012/T2	BL5	net939	I0/I3012/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2990/T2	BL5	net938	I0/I2990/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3003/T3	I0/I3003/net049	net946	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2993/T3	I0/I2993/net049	net945	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3019/T3	I0/I3019/net049	net944	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3013/T3	I0/I3013/net049	net943	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2999/T3	I0/I2999/net049	net942	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2992/T3	I0/I2992/net049	net941	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3015/T3	I0/I3015/net049	net940	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3012/T3	I0/I3012/net049	net939	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2990/T3	I0/I2990/net049	net938	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3035/T2	BL6	net946	I0/I3035/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3025/T2	BL6	net945	I0/I3025/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3051/T2	BL6	net944	I0/I3051/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3045/T2	BL6	net943	I0/I3045/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3031/T2	BL6	net942	I0/I3031/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3024/T2	BL6	net941	I0/I3024/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3047/T2	BL6	net940	I0/I3047/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3044/T2	BL6	net939	I0/I3044/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3022/T2	BL6	net938	I0/I3022/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3035/T5	I0/I3035/net13	I0/I3035/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3025/T5	I0/I3025/net13	I0/I3025/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3051/T5	I0/I3051/net13	I0/I3051/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3045/T5	I0/I3045/net13	I0/I3045/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3031/T5	I0/I3031/net13	I0/I3031/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3024/T5	I0/I3024/net13	I0/I3024/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3047/T5	I0/I3047/net13	I0/I3047/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3044/T5	I0/I3044/net13	I0/I3044/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3022/T5	I0/I3022/net13	I0/I3022/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3035/T4	vss	I0/I3035/net13	I0/I3035/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3025/T4	vss	I0/I3025/net13	I0/I3025/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3051/T4	vss	I0/I3051/net13	I0/I3051/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3045/T4	vss	I0/I3045/net13	I0/I3045/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3031/T4	vss	I0/I3031/net13	I0/I3031/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3024/T4	vss	I0/I3024/net13	I0/I3024/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3047/T4	vss	I0/I3047/net13	I0/I3047/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3044/T4	vss	I0/I3044/net13	I0/I3044/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3022/T4	vss	I0/I3022/net13	I0/I3022/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3035/T3	I0/I3035/net049	net946	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3025/T3	I0/I3025/net049	net945	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3051/T3	I0/I3051/net049	net944	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3045/T3	I0/I3045/net049	net943	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3031/T3	I0/I3031/net049	net942	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3024/T3	I0/I3024/net049	net941	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3047/T3	I0/I3047/net049	net940	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3044/T3	I0/I3044/net049	net939	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3022/T3	I0/I3022/net049	net938	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3067/T2	BL7	net946	I0/I3067/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3057/T2	BL7	net945	I0/I3057/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3083/T2	BL7	net944	I0/I3083/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3077/T2	BL7	net943	I0/I3077/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3063/T2	BL7	net942	I0/I3063/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3056/T2	BL7	net941	I0/I3056/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3079/T2	BL7	net940	I0/I3079/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3076/T2	BL7	net939	I0/I3076/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3054/T2	BL7	net938	I0/I3054/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T1	net955	I1/net1308	vss	vss	nfet	L=0.12U	W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.824e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2862/T5	I0/I2862/net13	I0/I2862/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2862/T2	BL1	net955	I0/I2862/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I84/T3	I0/I84/net049	net955	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I84/T4	vss	I0/I84/net13	I0/I84/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I84/T5	I0/I84/net13	I0/I84/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I84/T2	BL0	net955	I0/I84/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3068/T3	I0/I3068/net049	net955	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3068/T4	vss	I0/I3068/net13	I0/I3068/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3068/T5	I0/I3068/net13	I0/I3068/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2862/T4	vss	I0/I2862/net13	I0/I2862/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2926/T3	I0/I2926/net049	net955	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2926/T4	vss	I0/I2926/net13	I0/I2926/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2926/T5	I0/I2926/net13	I0/I2926/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2926/T2	BL3	net955	I0/I2926/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2894/T3	I0/I2894/net049	net955	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2894/T4	vss	I0/I2894/net13	I0/I2894/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2894/T5	I0/I2894/net13	I0/I2894/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2894/T2	BL2	net955	I0/I2894/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2862/T3	I0/I2862/net049	net955	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I82/T3	I0/I82/net049	net954	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I82/T4	vss	I0/I82/net13	I0/I82/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I82/T5	I0/I82/net13	I0/I82/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I82/T2	BL0	net954	I0/I82/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3060/T3	I0/I3060/net049	net954	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3060/T4	vss	I0/I3060/net13	I0/I3060/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3060/T5	I0/I3060/net13	I0/I3060/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2895/T4	vss	I0/I2895/net13	I0/I2895/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2895/T5	I0/I2895/net13	I0/I2895/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2895/T2	BL2	net954	I0/I2895/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2866/T3	I0/I2866/net049	net954	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2866/T4	vss	I0/I2866/net13	I0/I2866/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2866/T5	I0/I2866/net13	I0/I2866/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2866/T2	BL1	net954	I0/I2866/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2895/T3	I0/I2895/net049	net954	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T66	net954	I1/net1260	vss	vss	nfet	L=0.12U	W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2934/T3	I0/I2934/net049	net954	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2934/T4	vss	I0/I2934/net13	I0/I2934/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2934/T5	I0/I2934/net13	I0/I2934/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2934/T2	BL3	net954	I0/I2934/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T89	net953	I1/net1220	vss	vss	nfet	L=0.12U	W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.056e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2888/T5	I0/I2888/net13	I0/I2888/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2888/T2	BL1	net953	I0/I2888/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I6/T3	I0/I6/net049	net953	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I6/T4	vss	I0/I6/net13	I0/I6/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I6/T5	I0/I6/net13	I0/I6/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I6/T2	BL0	net953	I0/I6/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3059/T3	I0/I3059/net049	net953	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3059/T4	vss	I0/I3059/net13	I0/I3059/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3059/T5	I0/I3059/net13	I0/I3059/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2888/T4	vss	I0/I2888/net13	I0/I2888/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2933/T3	I0/I2933/net049	net953	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2933/T4	vss	I0/I2933/net13	I0/I2933/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2933/T5	I0/I2933/net13	I0/I2933/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2933/T2	BL3	net953	I0/I2933/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2909/T3	I0/I2909/net049	net953	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2909/T4	vss	I0/I2909/net13	I0/I2909/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2909/T5	I0/I2909/net13	I0/I2909/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2909/T2	BL2	net953	I0/I2909/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2888/T3	I0/I2888/net049	net953	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I5/T3	I0/I5/net049	net952	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I5/T4	vss	I0/I5/net13	I0/I5/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I5/T5	I0/I5/net13	I0/I5/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I5/T2	BL0	net952	I0/I5/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3084/T3	I0/I3084/net049	net952	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3084/T4	vss	I0/I3084/net13	I0/I3084/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3084/T5	I0/I3084/net13	I0/I3084/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2923/T4	vss	I0/I2923/net13	I0/I2923/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2923/T5	I0/I2923/net13	I0/I2923/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2923/T2	BL2	net952	I0/I2923/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2893/T3	I0/I2893/net049	net952	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2893/T4	vss	I0/I2893/net13	I0/I2893/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2893/T5	I0/I2893/net13	I0/I2893/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2893/T2	BL1	net952	I0/I2893/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2923/T3	I0/I2923/net049	net952	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T110	net952	I1/net1176	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2951/T3	I0/I2951/net049	net952	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2951/T4	vss	I0/I2951/net13	I0/I2951/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2951/T5	I0/I2951/net13	I0/I2951/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2951/T2	BL3	net952	I0/I2951/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T175	net951	I1/net1324	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=8.6e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3065/T3	I0/I3065/net049	net951	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3080/T3	I0/I3080/net049	net950	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3065/T4	vss	I0/I3065/net13	I0/I3065/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3080/T4	vss	I0/I3080/net13	I0/I3080/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3065/T5	I0/I3065/net13	I0/I3065/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3080/T5	I0/I3080/net13	I0/I3080/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3078/T3	I0/I3078/net049	net949	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3078/T4	vss	I0/I3078/net13	I0/I3078/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3078/T5	I0/I3078/net13	I0/I3078/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3074/T3	I0/I3074/net049	net948	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3066/T3	I0/I3066/net049	net947	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3074/T4	vss	I0/I3074/net13	I0/I3074/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3066/T4	vss	I0/I3066/net13	I0/I3066/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3074/T5	I0/I3074/net13	I0/I3074/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3066/T5	I0/I3066/net13	I0/I3066/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2821/T5	I0/I2821/net13	I0/I2821/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2812/T5	I0/I2812/net13	I0/I2812/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2825/T5	I0/I2825/net13	I0/I2825/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2805/T5	I0/I2805/net13	I0/I2805/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2826/T5	I0/I2826/net13	I0/I2826/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2821/T2	BL0	net951	I0/I2821/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2812/T2	BL0	net950	I0/I2812/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2825/T2	BL0	net949	I0/I2825/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2805/T2	BL0	net948	I0/I2805/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2826/T2	BL0	net947	I0/I2826/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2821/T3	I0/I2821/net049	net951	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2812/T3	I0/I2812/net049	net950	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2825/T3	I0/I2825/net049	net949	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2805/T3	I0/I2805/net049	net948	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2826/T3	I0/I2826/net049	net947	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2821/T4	vss	I0/I2821/net13	I0/I2821/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2812/T4	vss	I0/I2812/net13	I0/I2812/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2825/T4	vss	I0/I2825/net13	I0/I2825/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2805/T4	vss	I0/I2805/net13	I0/I2805/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2826/T4	vss	I0/I2826/net13	I0/I2826/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2871/T5	I0/I2871/net13	I0/I2871/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2877/T5	I0/I2877/net13	I0/I2877/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2879/T5	I0/I2879/net13	I0/I2879/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2886/T5	I0/I2886/net13	I0/I2886/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2872/T5	I0/I2872/net13	I0/I2872/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2871/T2	BL1	net951	I0/I2871/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2877/T2	BL1	net950	I0/I2877/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2879/T2	BL1	net949	I0/I2879/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2886/T2	BL1	net948	I0/I2886/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2872/T2	BL1	net947	I0/I2872/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2871/T3	I0/I2871/net049	net951	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2877/T3	I0/I2877/net049	net950	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2879/T3	I0/I2879/net049	net949	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2886/T3	I0/I2886/net049	net948	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2872/T3	I0/I2872/net049	net947	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2871/T4	vss	I0/I2871/net13	I0/I2871/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2877/T4	vss	I0/I2877/net13	I0/I2877/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2879/T4	vss	I0/I2879/net13	I0/I2879/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2886/T4	vss	I0/I2886/net13	I0/I2886/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2872/T4	vss	I0/I2872/net13	I0/I2872/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2903/T4	vss	I0/I2903/net13	I0/I2903/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2922/T4	vss	I0/I2922/net13	I0/I2922/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2903/T5	I0/I2903/net13	I0/I2903/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2922/T5	I0/I2922/net13	I0/I2922/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2903/T2	BL2	net951	I0/I2903/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2922/T2	BL2	net950	I0/I2922/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2919/T4	vss	I0/I2919/net13	I0/I2919/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2919/T5	I0/I2919/net13	I0/I2919/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2919/T2	BL2	net949	I0/I2919/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2910/T4	vss	I0/I2910/net13	I0/I2910/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2905/T4	vss	I0/I2905/net13	I0/I2905/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2910/T5	I0/I2910/net13	I0/I2910/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2905/T5	I0/I2905/net13	I0/I2905/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2910/T2	BL2	net948	I0/I2910/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2905/T2	BL2	net947	I0/I2905/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2903/T3	I0/I2903/net049	net951	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2922/T3	I0/I2922/net049	net950	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2919/T3	I0/I2919/net049	net949	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2910/T3	I0/I2910/net049	net948	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2905/T3	I0/I2905/net049	net947	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2940/T5	I0/I2940/net13	I0/I2940/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2956/T5	I0/I2956/net13	I0/I2956/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2957/T5	I0/I2957/net13	I0/I2957/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2936/T5	I0/I2936/net13	I0/I2936/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2941/T5	I0/I2941/net13	I0/I2941/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2940/T2	BL3	net951	I0/I2940/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2956/T2	BL3	net950	I0/I2956/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2957/T2	BL3	net949	I0/I2957/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2936/T2	BL3	net948	I0/I2936/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2941/T2	BL3	net947	I0/I2941/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2940/T3	I0/I2940/net049	net951	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2956/T3	I0/I2956/net049	net950	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2957/T3	I0/I2957/net049	net949	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2936/T3	I0/I2936/net049	net948	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2941/T3	I0/I2941/net049	net947	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2940/T4	vss	I0/I2940/net13	I0/I2940/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2956/T4	vss	I0/I2956/net13	I0/I2956/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2957/T4	vss	I0/I2957/net13	I0/I2957/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2936/T4	vss	I0/I2936/net13	I0/I2936/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2941/T4	vss	I0/I2941/net13	I0/I2941/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T185	net950	I1/net1492	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.032e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T192	net949	I1/net1436	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T205	net948	I1/net1452	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T270	net947	I1/net1644	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3067/T3	I0/I3067/net049	net946	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3057/T3	I0/I3057/net049	net945	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3067/T4	vss	I0/I3067/net13	I0/I3067/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3057/T4	vss	I0/I3057/net13	I0/I3057/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3067/T5	I0/I3067/net13	I0/I3067/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3057/T5	I0/I3057/net13	I0/I3057/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3083/T3	I0/I3083/net049	net944	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3083/T4	vss	I0/I3083/net13	I0/I3083/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3083/T5	I0/I3083/net13	I0/I3083/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3077/T3	I0/I3077/net049	net943	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3063/T3	I0/I3063/net049	net942	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3077/T4	vss	I0/I3077/net13	I0/I3077/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3063/T4	vss	I0/I3063/net13	I0/I3063/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3077/T5	I0/I3077/net13	I0/I3077/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3063/T5	I0/I3063/net13	I0/I3063/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2816/T5	I0/I2816/net13	I0/I2816/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2803/T5	I0/I2803/net13	I0/I2803/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2811/T5	I0/I2811/net13	I0/I2811/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2813/T5	I0/I2813/net13	I0/I2813/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2827/T5	I0/I2827/net13	I0/I2827/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2816/T2	BL0	net946	I0/I2816/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2803/T2	BL0	net945	I0/I2803/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2811/T2	BL0	net944	I0/I2811/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2813/T2	BL0	net943	I0/I2813/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2827/T2	BL0	net942	I0/I2827/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2816/T3	I0/I2816/net049	net946	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2803/T3	I0/I2803/net049	net945	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2811/T3	I0/I2811/net049	net944	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2813/T3	I0/I2813/net049	net943	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2827/T3	I0/I2827/net049	net942	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2816/T4	vss	I0/I2816/net13	I0/I2816/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2803/T4	vss	I0/I2803/net13	I0/I2803/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2811/T4	vss	I0/I2811/net13	I0/I2811/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2813/T4	vss	I0/I2813/net13	I0/I2813/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2827/T4	vss	I0/I2827/net13	I0/I2827/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2887/T5	I0/I2887/net13	I0/I2887/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2889/T5	I0/I2889/net13	I0/I2889/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2880/T5	I0/I2880/net13	I0/I2880/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2881/T5	I0/I2881/net13	I0/I2881/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2865/T5	I0/I2865/net13	I0/I2865/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2887/T2	BL1	net946	I0/I2887/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2889/T2	BL1	net945	I0/I2889/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2880/T2	BL1	net944	I0/I2880/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2881/T2	BL1	net943	I0/I2881/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2865/T2	BL1	net942	I0/I2865/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2887/T3	I0/I2887/net049	net946	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2889/T3	I0/I2889/net049	net945	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2880/T3	I0/I2880/net049	net944	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2881/T3	I0/I2881/net049	net943	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2865/T3	I0/I2865/net049	net942	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2887/T4	vss	I0/I2887/net13	I0/I2887/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2889/T4	vss	I0/I2889/net13	I0/I2889/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2880/T4	vss	I0/I2880/net13	I0/I2880/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2881/T4	vss	I0/I2881/net13	I0/I2881/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2865/T4	vss	I0/I2865/net13	I0/I2865/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2920/T4	vss	I0/I2920/net13	I0/I2920/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2915/T4	vss	I0/I2915/net13	I0/I2915/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2920/T5	I0/I2920/net13	I0/I2920/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2915/T5	I0/I2915/net13	I0/I2915/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2920/T2	BL2	net946	I0/I2920/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2915/T2	BL2	net945	I0/I2915/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2902/T4	vss	I0/I2902/net13	I0/I2902/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2902/T5	I0/I2902/net13	I0/I2902/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2902/T2	BL2	net944	I0/I2902/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2901/T4	vss	I0/I2901/net13	I0/I2901/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2914/T4	vss	I0/I2914/net13	I0/I2914/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2901/T5	I0/I2901/net13	I0/I2901/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2914/T5	I0/I2914/net13	I0/I2914/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2901/T2	BL2	net943	I0/I2901/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2914/T2	BL2	net942	I0/I2914/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2920/T3	I0/I2920/net049	net946	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2915/T3	I0/I2915/net049	net945	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2902/T3	I0/I2902/net049	net944	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2901/T3	I0/I2901/net049	net943	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2914/T3	I0/I2914/net049	net942	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2953/T5	I0/I2953/net13	I0/I2953/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2949/T5	I0/I2949/net13	I0/I2949/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2938/T5	I0/I2938/net13	I0/I2938/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2935/T5	I0/I2935/net13	I0/I2935/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2947/T5	I0/I2947/net13	I0/I2947/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2953/T2	BL3	net946	I0/I2953/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2949/T2	BL3	net945	I0/I2949/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2938/T2	BL3	net944	I0/I2938/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2935/T2	BL3	net943	I0/I2935/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2947/T2	BL3	net942	I0/I2947/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2953/T3	I0/I2953/net049	net946	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2949/T3	I0/I2949/net049	net945	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2938/T3	I0/I2938/net049	net944	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2935/T3	I0/I2935/net049	net943	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2947/T3	I0/I2947/net049	net942	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2953/T4	vss	I0/I2953/net13	I0/I2953/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2949/T4	vss	I0/I2949/net13	I0/I2949/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2938/T4	vss	I0/I2938/net13	I0/I2938/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2935/T4	vss	I0/I2935/net13	I0/I2935/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2947/T4	vss	I0/I2947/net13	I0/I2947/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T260	net946	I1/net1616	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T253	net945	I1/net1588	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T240	net944	I1/net1544	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T303	net943	I1/net1672	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T313	net942	I1/net1464	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2890/T5	I0/I2890/net13	I0/I2890/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2890/T2	BL1	net941	I0/I2890/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2804/T3	I0/I2804/net049	net941	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2804/T4	vss	I0/I2804/net13	I0/I2804/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2804/T5	I0/I2804/net13	I0/I2804/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2804/T2	BL0	net941	I0/I2804/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3056/T3	I0/I3056/net049	net941	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3056/T4	vss	I0/I3056/net13	I0/I3056/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3056/T5	I0/I3056/net13	I0/I3056/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2890/T4	vss	I0/I2890/net13	I0/I2890/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2950/T3	I0/I2950/net049	net941	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2950/T4	vss	I0/I2950/net13	I0/I2950/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2950/T5	I0/I2950/net13	I0/I2950/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2950/T2	BL3	net941	I0/I2950/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2913/T3	I0/I2913/net049	net941	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2913/T4	vss	I0/I2913/net13	I0/I2913/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2913/T5	I0/I2913/net13	I0/I2913/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2913/T2	BL2	net941	I0/I2913/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2890/T3	I0/I2890/net049	net941	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T320	net941	I1/net1816	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2891/T5	I0/I2891/net13	I0/I2891/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2891/T2	BL1	net940	I0/I2891/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2802/T3	I0/I2802/net049	net940	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2802/T4	vss	I0/I2802/net13	I0/I2802/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2802/T5	I0/I2802/net13	I0/I2802/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2802/T2	BL0	net940	I0/I2802/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3079/T3	I0/I3079/net049	net940	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3079/T4	vss	I0/I3079/net13	I0/I3079/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3079/T5	I0/I3079/net13	I0/I3079/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2891/T4	vss	I0/I2891/net13	I0/I2891/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2943/T3	I0/I2943/net049	net940	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2943/T4	vss	I0/I2943/net13	I0/I2943/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2943/T5	I0/I2943/net13	I0/I2943/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2943/T2	BL3	net940	I0/I2943/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2908/T3	I0/I2908/net049	net940	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2908/T4	vss	I0/I2908/net13	I0/I2908/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2908/T5	I0/I2908/net13	I0/I2908/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2908/T2	BL2	net940	I0/I2908/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2891/T3	I0/I2891/net049	net940	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T333	net940	I1/net1852	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3076/T3	I0/I3076/net049	net939	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3054/T3	I0/I3054/net049	net938	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3076/T4	vss	I0/I3076/net13	I0/I3076/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3054/T4	vss	I0/I3054/net13	I0/I3054/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3076/T5	I0/I3076/net13	I0/I3076/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3054/T5	I0/I3054/net13	I0/I3054/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2820/T3	I0/I2820/net049	net939	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2800/T3	I0/I2800/net049	net938	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2820/T4	vss	I0/I2820/net13	I0/I2820/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2800/T4	vss	I0/I2800/net13	I0/I2800/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2820/T5	I0/I2820/net13	I0/I2820/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2800/T5	I0/I2800/net13	I0/I2800/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2820/T2	BL0	net939	I0/I2820/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2800/T2	BL0	net938	I0/I2800/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2875/T3	I0/I2875/net049	net939	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2883/T3	I0/I2883/net049	net938	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2875/T4	vss	I0/I2875/net13	I0/I2875/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2883/T4	vss	I0/I2883/net13	I0/I2883/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2875/T5	I0/I2875/net13	I0/I2875/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2883/T5	I0/I2883/net13	I0/I2883/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2875/T2	BL1	net939	I0/I2875/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2883/T2	BL1	net938	I0/I2883/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2912/T4	vss	I0/I2912/net13	I0/I2912/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2918/T4	vss	I0/I2918/net13	I0/I2918/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2912/T5	I0/I2912/net13	I0/I2912/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2918/T5	I0/I2918/net13	I0/I2918/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2912/T2	BL2	net939	I0/I2912/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2918/T2	BL2	net938	I0/I2918/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2912/T3	I0/I2912/net049	net939	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2918/T3	I0/I2918/net049	net938	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T398	net939	I1/net1904	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T388	net938	I1/net1772	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2948/T3	I0/I2948/net049	net939	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2952/T3	I0/I2952/net049	net938	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2948/T4	vss	I0/I2948/net13	I0/I2948/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2952/T4	vss	I0/I2952/net13	I0/I2952/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2948/T5	I0/I2948/net13	I0/I2948/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2952/T5	I0/I2952/net13	I0/I2952/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2948/T2	BL3	net939	I0/I2948/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2952/T2	BL3	net938	I0/I2952/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI159/T7	vss	I159/net28	clkout	vss	nfet	L=0.12U
+ W=17.29U
+ AD=5.5328P	AS=5.5328P	PD=35.22U	PS=35.22U
+ wt=1.729e-05 wf=1.729e-05 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.0988e-12 panw6=9.6e-15 panw10=7.2e-14 nrs=0.0127573 nrd=0.0127573 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T8	I1/net1292	I1/net160	I1/net168	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=9.24e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T9	I1/net168	I1/a3bar	I1/net164	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=6.51e-14 panw8=2.4e-14 panw7=1.92e-14 panw10=2.85e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T10	I1/net164	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 panw10=6.84e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T63	I1/net1248	I1/net160	I1/net108	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T7	I1/net176	I1/net1292	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=6.72e-14 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI159/T6	vss	I159/net32	I159/net28	vss	nfet	L=0.12U
+ W=4.6U
+ AD=1.472P	AS=1.472P	PD=9.84U	PS=9.84U
+ wt=4.6e-06 wf=4.6e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.76e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0482986 nrd=0.0482986 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T2	I1/net1308	I1/net176	I1/net180	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=3.204e-13 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T3	I1/net180	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.209e-13 panw8=2.4e-14 panw7=2.16e-14 panw10=1.955e-13 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T65	I1/net1260	I1/net112	I1/net132	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T60	I1/net112	I1/net1248	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T95	I1/net76	I1/net1208	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T104	I1/net72	I1/net1188	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T64	I1/net132	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T90	I1/net1220	I1/net76	I1/net92	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T91	I1/net92	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T109	I1/net1176	I1/net72	I1/net56	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T108	I1/net56	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T62	I1/net108	I1/a3bar	I1/net104	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T61	I1/net104	I1/a4	vss	vss	nfet	L=0.12U	W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T92	I1/net1208	I1/net160	I1/net84	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T93	I1/net84	I1/a3	I1/net80	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T94	I1/net80	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T107	I1/net1188	I1/net160	I1/net64	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T106	I1/net64	I1/a3	I1/net68	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T105	I1/net68	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T178	I1/net412	I1/net1420	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T189	I1/net284	I1/net1328	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T176	I1/net1324	I1/net412	I1/net324	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T177	I1/net324	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T186	I1/net1492	I1/net284	I1/net200	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T187	I1/net200	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T193	I1/net1436	I1/net420	I1/net304	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T198	I1/net420	I1/net1496	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T199	I1/net352	I1/net1488	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T194	I1/net304	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T204	I1/net1452	I1/net352	I1/net400	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T203	I1/net400	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T269	I1/net1644	I1/net532	I1/net536	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T179	I1/net1420	I1/net316	I1/net396	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T180	I1/net396	I1/a3bar	I1/net380	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T181	I1/net380	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T188	I1/net1328	I1/net316	I1/net364	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T190	I1/net364	I1/a3bar	I1/net252	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T191	I1/net252	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T195	I1/net1496	I1/net316	I1/net368	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T196	I1/net368	I1/a3	I1/net384	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T197	I1/net384	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T202	I1/net1488	I1/net316	I1/net340	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T201	I1/net340	I1/a3	I1/net360	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T200	I1/net360	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T266	I1/net1628	I1/net516	I1/net524	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T267	I1/net532	I1/net1628	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T256	I1/net492	I1/net1604	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T247	I1/net456	I1/net1576	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T268	I1/net536	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T259	I1/net1616	I1/net492	I1/net500	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T258	I1/net500	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T252	I1/net1588	I1/net456	I1/net472	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T251	I1/net472	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T246	I1/net452	I1/net1556	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T306	I1/net600	I1/net1840	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T241	I1/net1544	I1/net452	I1/net436	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T242	I1/net436	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T304	I1/net1672	I1/net600	I1/net724	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T305	I1/net724	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T317	I1/net768	I1/net1792	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T326	I1/net704	I1/net1352	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T314	I1/net1464	I1/net768	I1/net772	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T315	I1/net772	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T321	I1/net1816	I1/net704	I1/net688	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T322	I1/net688	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T332	I1/net1852	I1/net708	I1/net344	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T327	I1/net708	I1/net1880	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T395	I1/net788	I1/net1716	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T384	I1/net796	I1/net1800	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T331	I1/net344	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T397	I1/net1904	I1/net788	I1/net628	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T396	I1/net628	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T387	I1/net1772	I1/net796	I1/net632	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T386	I1/net632	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T265	I1/net524	I1/a3bar	I1/net520	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T264	I1/net520	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T257	I1/net1604	I1/net516	I1/net488	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T255	I1/net488	I1/a3bar	I1/net484	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T254	I1/net484	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T250	I1/net1576	I1/net516	I1/net464	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T249	I1/net464	I1/a3	I1/net460	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T248	I1/net460	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T243	I1/net1556	I1/net516	I1/net444	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T244	I1/net444	I1/a3	I1/net448	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T245	I1/net448	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T307	I1/net1840	I1/net776	I1/net604	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T308	I1/net604	I1/a3bar	I1/net784	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T309	I1/net784	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T316	I1/net1792	I1/net776	I1/net680	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T318	I1/net680	I1/a3bar	I1/net672	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T319	I1/net672	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T323	I1/net1352	I1/net776	I1/net692	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T324	I1/net692	I1/a3	I1/net696	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T325	I1/net696	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T330	I1/net1880	I1/net776	I1/net564	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T329	I1/net564	I1/a3	I1/net568	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T328	I1/net568	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T394	I1/net1716	I1/net616	I1/net736	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T393	I1/net736	I1/a3bar	I1/net624	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T392	I1/net624	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T385	I1/net1800	I1/net616	I1/net792	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T383	I1/net792	I1/a3bar	I1/net808	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T382	I1/net808	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T18	I1/net148	I1/a2bar	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T184	I1/net388	I1/a2	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T17	I1/net152	I1/a1bar	I1/net148	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T183	I1/net376	I1/a1bar	I1/net388	vss	nfet
+ L=0.12U	W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T15	I1/net160	I1/net1284	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T182	I1/net316	I1/net1460	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T16	I1/net1284	I1/a0bar	I1/net152	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T206	I1/net1460	I1/a0bar	I1/net376	vss	nfet
+ L=0.12U	W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T263	I1/net516	I1/net1656	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T261	I1/net296	I1/a2bar	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T312	I1/net584	I1/a2	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T262	I1/net512	I1/a1	I1/net296	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T311	I1/net780	I1/a1	I1/net584	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T310	I1/net776	I1/net1820	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T391	I1/net616	I1/net1860	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T239	I1/net1656	I1/a0bar	I1/net512	vss	nfet
+ L=0.12U	W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T334	I1/net1820	I1/a0bar	I1/net780	vss	nfet
+ L=0.12U	W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T31	vss	addr0	I1/a0bar	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T32	vss	addr1	I1/a1bar	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T25	I1/net156	addr0	vss	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1188P	AS=0.1221P	PD=1.38U	PS=1.4U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T48	I1/net144	addr1	vss	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1188P	AS=0.1221P	PD=1.38U	PS=1.4U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI159/T4	vss	clk	I159/net36	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=4.32e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T24	I1/a0	I1/net156	vss	vss	nfet	L=0.12U	W=0.57U
+ AD=0.2052P	AS=0.2109P	PD=1.86U	PS=1.88U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T26	I1/a1	I1/net144	vss	vss	nfet	L=0.12U	W=0.57U
+ AD=0.2052P	AS=0.2109P	PD=1.86U	PS=1.88U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI159/T5	vss	I159/net36	I159/net32	vss	nfet	L=0.12U
+ W=1.24U
+ AD=0.3968P	AS=0.3968P	PD=3.12U	PS=3.12U
+ wt=1.24e-06 wf=1.24e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.76e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=4.1e-14 nrs=0.1841 nrd=0.1841 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T45	vss	I1/net264	I1/net260	vss	nfet	L=0.12U
+ W=0.83U
+ AD=0.3071P	AS=0.2988P	PD=2.4U	PS=2.38U
+ wt=8.3e-07 wf=8.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.56e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=9.96e-14 nrs=0.280255 nrd=0.280255 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T43	I1/net264	I1/net124	vss	vss	nfet	L=0.12U
+ W=0.52U
+ AD=0.1872P	AS=0.1924P	PD=1.76U	PS=1.78U
+ wt=5.2e-07 wf=5.2e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.6e-14 nrs=0.463158 nrd=0.463158 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T33	vss	addr2	I1/a2bar	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T55	I1/net116	addr2	vss	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1188P	AS=0.1221P	PD=1.38U	PS=1.4U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T29	I1/a2	I1/net116	vss	vss	nfet	L=0.12U	W=0.57U
+ AD=0.2052P	AS=0.2109P	PD=1.86U	PS=1.88U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T54	I1/a3	I1/net260	vss	vss	nfet	L=0.12U	W=2.05U
+ AD=0.738P	AS=0.7585P	PD=4.82U	PS=4.84U
+ wt=2.05e-06 wf=2.05e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.916e-13 nrs=0.109726 nrd=0.109726 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T34	vss	addr3	I1/net124	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T69	vss	addr3	I1/net328	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.96e-14 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T46	vss	I1/net212	I1/net256	vss	nfet	L=0.12U
+ W=0.83U
+ AD=0.3071P	AS=0.2988P	PD=2.4U	PS=2.38U
+ wt=8.3e-07 wf=8.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.56e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=9.96e-14 nrs=0.280255 nrd=0.280255 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T41	vss	addr4	I1/net120	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T96	vss	addr4	I1/net216	vss	nfet	L=0.12U	W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.96e-14 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T67	I1/net320	I1/net328	vss	vss	nfet	L=0.12U
+ W=0.83U
+ AD=0.2988P	AS=0.3071P	PD=2.38U	PS=2.4U
+ wt=8.3e-07 wf=8.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-15 panw8=3e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.48e-14 nrs=0.280255 nrd=0.280255 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T44	I1/net212	I1/net120	vss	vss	nfet	L=0.12U
+ W=0.52U
+ AD=0.1872P	AS=0.1924P	PD=1.76U	PS=1.78U
+ wt=5.2e-07 wf=5.2e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.6e-14 nrs=0.463158 nrd=0.463158 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T59	I1/a3bar	I1/net320	vss	vss	nfet	L=0.12U
+ W=2.05U
+ AD=0.738P	AS=0.7585P	PD=4.82U	PS=4.84U
+ wt=2.05e-06 wf=2.05e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.296e-13 nrs=0.109726 nrd=0.109726 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T56	I1/a4	I1/net256	vss	vss	nfet	L=0.12U	W=2.05U
+ AD=0.738P	AS=0.7585P	PD=4.82U	PS=4.84U
+ wt=2.05e-06 wf=2.05e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.916e-13 nrs=0.109726 nrd=0.109726 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T88	I1/a4bar	I1/net336	vss	vss	nfet	L=0.12U
+ W=2.05U
+ AD=0.738P	AS=0.7585P	PD=4.82U	PS=4.84U
+ wt=2.05e-06 wf=2.05e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.296e-13 nrs=0.109726 nrd=0.109726 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T87	I1/net336	I1/net216	vss	vss	nfet	L=0.12U
+ W=0.83U
+ AD=0.2988P	AS=0.3071P	PD=2.38U	PS=2.4U
+ wt=8.3e-07 wf=8.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.56e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.48e-14 nrs=0.280255 nrd=0.280255 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3151/T3	I0/I3151/net049	net937	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3151/T4	vss	I0/I3151/net13	I0/I3151/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3151/T5	I0/I3151/net13	I0/I3151/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3151/T2	BL10	net937	I0/I3151/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3119/T3	I0/I3119/net049	net937	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3119/T4	vss	I0/I3119/net13	I0/I3119/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3119/T5	I0/I3119/net13	I0/I3119/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3119/T2	BL9	net937	I0/I3119/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3087/T3	I0/I3087/net049	net937	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3087/T4	vss	I0/I3087/net13	I0/I3087/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3087/T5	I0/I3087/net13	I0/I3087/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3158/T3	I0/I3158/net049	net936	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3158/T4	vss	I0/I3158/net13	I0/I3158/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3158/T5	I0/I3158/net13	I0/I3158/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3158/T2	BL10	net936	I0/I3158/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3126/T3	I0/I3126/net049	net936	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3126/T4	vss	I0/I3126/net13	I0/I3126/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3126/T5	I0/I3126/net13	I0/I3126/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3126/T2	BL9	net936	I0/I3126/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3094/T3	I0/I3094/net049	net936	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3094/T4	vss	I0/I3094/net13	I0/I3094/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3094/T5	I0/I3094/net13	I0/I3094/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I120/T5	I0/I120/net13	I0/I120/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I120/T2	BL4	net937	I0/I120/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3183/T3	I0/I3183/net049	net937	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3183/T4	vss	I0/I3183/net13	I0/I3183/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3183/T5	I0/I3183/net13	I0/I3183/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3183/T2	BL11	net937	I0/I3183/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I113/T5	I0/I113/net13	I0/I113/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I113/T2	BL4	net936	I0/I113/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3190/T3	I0/I3190/net049	net936	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3190/T4	vss	I0/I3190/net13	I0/I3190/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3190/T5	I0/I3190/net13	I0/I3190/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3190/T2	BL11	net936	I0/I3190/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2991/T3	I0/I2991/net049	net937	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2991/T4	vss	I0/I2991/net13	I0/I2991/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2991/T5	I0/I2991/net13	I0/I2991/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2991/T2	BL5	net937	I0/I2991/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I120/T3	I0/I120/net049	net937	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I120/T4	vss	I0/I120/net13	I0/I120/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2998/T3	I0/I2998/net049	net936	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2998/T4	vss	I0/I2998/net13	I0/I2998/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2998/T5	I0/I2998/net13	I0/I2998/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2998/T2	BL5	net936	I0/I2998/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I113/T3	I0/I113/net049	net936	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I113/T4	vss	I0/I113/net13	I0/I113/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3055/T5	I0/I3055/net13	I0/I3055/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3055/T2	BL7	net937	I0/I3055/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3023/T3	I0/I3023/net049	net937	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3023/T4	vss	I0/I3023/net13	I0/I3023/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3023/T5	I0/I3023/net13	I0/I3023/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3023/T2	BL6	net937	I0/I3023/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3062/T5	I0/I3062/net13	I0/I3062/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3062/T2	BL7	net936	I0/I3062/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3030/T3	I0/I3030/net049	net936	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3030/T4	vss	I0/I3030/net13	I0/I3030/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3030/T5	I0/I3030/net13	I0/I3030/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3030/T2	BL6	net936	I0/I3030/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2810/T3	I0/I2810/net049	net937	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2810/T4	vss	I0/I2810/net13	I0/I2810/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2810/T5	I0/I2810/net13	I0/I2810/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2810/T2	BL0	net937	I0/I2810/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3055/T3	I0/I3055/net049	net937	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3055/T4	vss	I0/I3055/net13	I0/I3055/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2809/T3	I0/I2809/net049	net936	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2809/T4	vss	I0/I2809/net13	I0/I2809/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2809/T5	I0/I2809/net13	I0/I2809/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2809/T2	BL0	net936	I0/I2809/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3062/T3	I0/I3062/net049	net936	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3062/T4	vss	I0/I3062/net13	I0/I3062/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2906/T5	I0/I2906/net13	I0/I2906/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2906/T2	BL2	net937	I0/I2906/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2885/T3	I0/I2885/net049	net937	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2885/T4	vss	I0/I2885/net13	I0/I2885/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2885/T5	I0/I2885/net13	I0/I2885/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2885/T2	BL1	net937	I0/I2885/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2916/T5	I0/I2916/net13	I0/I2916/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2916/T2	BL2	net936	I0/I2916/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2864/T3	I0/I2864/net049	net936	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2864/T4	vss	I0/I2864/net13	I0/I2864/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2864/T5	I0/I2864/net13	I0/I2864/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2864/T2	BL1	net936	I0/I2864/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2942/T3	I0/I2942/net049	net937	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2942/T4	vss	I0/I2942/net13	I0/I2942/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2942/T5	I0/I2942/net13	I0/I2942/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2942/T2	BL3	net937	I0/I2942/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2906/T3	I0/I2906/net049	net937	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2906/T4	vss	I0/I2906/net13	I0/I2906/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2932/T3	I0/I2932/net049	net936	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2932/T4	vss	I0/I2932/net13	I0/I2932/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2932/T5	I0/I2932/net13	I0/I2932/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2932/T2	BL3	net936	I0/I2932/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2916/T3	I0/I2916/net049	net936	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2916/T4	vss	I0/I2916/net13	I0/I2916/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T389	I1/net832	I1/a2bar	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T390	I1/net620	I1/a1bar	I1/net832	vss	nfet
+ L=0.12U	W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T367	I1/net1860	I1/a0	I1/net620	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T378	I1/net1780	I1/net616	I1/net660	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T377	I1/net660	I1/a3	I1/net652	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T376	I1/net652	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T375	I1/net732	I1/net1780	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T380	I1/net1752	I1/net732	I1/net740	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T379	I1/net740	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T381	net937	I1/net1752	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T97	vss	addr_en	I1/net02041	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1221P	AS=0.1188P	PD=1.4U	PS=1.38U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.96e-14 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T371	I1/net1484	I1/net616	I1/net204	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T372	I1/net204	I1/a3	I1/net608	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T373	I1/net608	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T374	I1/net812	I1/net1484	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T369	I1/net1708	I1/net812	I1/net196	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T370	I1/net196	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T368	net936	I1/net1708	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3160/T3	I0/I3160/net049	net935	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3160/T4	vss	I0/I3160/net13	I0/I3160/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3160/T5	I0/I3160/net13	I0/I3160/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3160/T2	BL10	net935	I0/I3160/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3128/T3	I0/I3128/net049	net935	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3128/T4	vss	I0/I3128/net13	I0/I3128/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3128/T5	I0/I3128/net13	I0/I3128/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3128/T2	BL9	net935	I0/I3128/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3096/T3	I0/I3096/net049	net935	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3096/T4	vss	I0/I3096/net13	I0/I3096/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3096/T5	I0/I3096/net13	I0/I3096/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I111/T5	I0/I111/net13	I0/I111/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I111/T2	BL4	net935	I0/I111/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3192/T3	I0/I3192/net049	net935	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3192/T4	vss	I0/I3192/net13	I0/I3192/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3192/T5	I0/I3192/net13	I0/I3192/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3192/T2	BL11	net935	I0/I3192/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3000/T3	I0/I3000/net049	net935	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3000/T4	vss	I0/I3000/net13	I0/I3000/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3000/T5	I0/I3000/net13	I0/I3000/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3000/T2	BL5	net935	I0/I3000/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I111/T3	I0/I111/net049	net935	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I111/T4	vss	I0/I111/net13	I0/I111/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3064/T5	I0/I3064/net13	I0/I3064/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3064/T2	BL7	net935	I0/I3064/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3032/T3	I0/I3032/net049	net935	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3032/T4	vss	I0/I3032/net13	I0/I3032/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3032/T5	I0/I3032/net13	I0/I3032/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3032/T2	BL6	net935	I0/I3032/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2801/T3	I0/I2801/net049	net935	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2801/T4	vss	I0/I2801/net13	I0/I2801/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2801/T5	I0/I2801/net13	I0/I2801/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2801/T2	BL0	net935	I0/I2801/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3064/T3	I0/I3064/net049	net935	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3064/T4	vss	I0/I3064/net13	I0/I3064/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2896/T5	I0/I2896/net13	I0/I2896/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2896/T2	BL2	net935	I0/I2896/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2867/T3	I0/I2867/net049	net935	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2867/T4	vss	I0/I2867/net13	I0/I2867/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2867/T5	I0/I2867/net13	I0/I2867/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2867/T2	BL1	net935	I0/I2867/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2928/T3	I0/I2928/net049	net935	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2928/T4	vss	I0/I2928/net13	I0/I2928/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2928/T5	I0/I2928/net13	I0/I2928/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2928/T2	BL3	net935	I0/I2928/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2896/T3	I0/I2896/net049	net935	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2896/T4	vss	I0/I2896/net13	I0/I2896/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T98	I1/net02030	I1/net02041	vss	vss	nfet	L=0.12U
+ W=1.18U
+ AD=0.4248P	AS=0.4366P	PD=3.08U	PS=3.1U
+ wt=1.18e-06 wf=1.18e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.512e-13 nrs=0.193833 nrd=0.193833 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T435	I1/net1960	I1/net880	I1/net872	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T432	I1/net1944	I1/net864	I1/net860	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3166/T3	I0/I3166/net049	net934	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3166/T4	vss	I0/I3166/net13	I0/I3166/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3166/T5	I0/I3166/net13	I0/I3166/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3166/T2	BL10	net934	I0/I3166/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3134/T3	I0/I3134/net049	net934	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3134/T4	vss	I0/I3134/net13	I0/I3134/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3134/T5	I0/I3134/net13	I0/I3134/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3134/T2	BL9	net934	I0/I3134/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3102/T3	I0/I3102/net049	net934	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3102/T4	vss	I0/I3102/net13	I0/I3102/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3102/T5	I0/I3102/net13	I0/I3102/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3168/T3	I0/I3168/net049	net933	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3168/T4	vss	I0/I3168/net13	I0/I3168/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3168/T5	I0/I3168/net13	I0/I3168/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3168/T2	BL10	net933	I0/I3168/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3136/T3	I0/I3136/net049	net933	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3136/T4	vss	I0/I3136/net13	I0/I3136/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3136/T5	I0/I3136/net13	I0/I3136/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3136/T2	BL9	net933	I0/I3136/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3104/T3	I0/I3104/net049	net933	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3104/T4	vss	I0/I3104/net13	I0/I3104/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3104/T5	I0/I3104/net13	I0/I3104/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3157/T3	I0/I3157/net049	net932	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3157/T4	vss	I0/I3157/net13	I0/I3157/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3157/T5	I0/I3157/net13	I0/I3157/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3157/T2	BL10	net932	I0/I3157/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3125/T3	I0/I3125/net049	net932	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3125/T4	vss	I0/I3125/net13	I0/I3125/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3125/T5	I0/I3125/net13	I0/I3125/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3125/T2	BL9	net932	I0/I3125/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3093/T3	I0/I3093/net049	net932	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3093/T4	vss	I0/I3093/net13	I0/I3093/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3093/T5	I0/I3093/net13	I0/I3093/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I105/T5	I0/I105/net13	I0/I105/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I105/T2	BL4	net934	I0/I105/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3198/T3	I0/I3198/net049	net934	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3198/T4	vss	I0/I3198/net13	I0/I3198/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3198/T5	I0/I3198/net13	I0/I3198/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3198/T2	BL11	net934	I0/I3198/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I103/T5	I0/I103/net13	I0/I103/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I103/T2	BL4	net933	I0/I103/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3200/T3	I0/I3200/net049	net933	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3200/T4	vss	I0/I3200/net13	I0/I3200/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3200/T5	I0/I3200/net13	I0/I3200/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3200/T2	BL11	net933	I0/I3200/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I114/T5	I0/I114/net13	I0/I114/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I114/T2	BL4	net932	I0/I114/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3189/T3	I0/I3189/net049	net932	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3189/T4	vss	I0/I3189/net13	I0/I3189/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3189/T5	I0/I3189/net13	I0/I3189/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3189/T2	BL11	net932	I0/I3189/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3006/T3	I0/I3006/net049	net934	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3006/T4	vss	I0/I3006/net13	I0/I3006/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3006/T5	I0/I3006/net13	I0/I3006/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3006/T2	BL5	net934	I0/I3006/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I105/T3	I0/I105/net049	net934	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I105/T4	vss	I0/I105/net13	I0/I105/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3008/T3	I0/I3008/net049	net933	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3008/T4	vss	I0/I3008/net13	I0/I3008/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3008/T5	I0/I3008/net13	I0/I3008/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3008/T2	BL5	net933	I0/I3008/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I103/T3	I0/I103/net049	net933	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I103/T4	vss	I0/I103/net13	I0/I103/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2997/T3	I0/I2997/net049	net932	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2997/T4	vss	I0/I2997/net13	I0/I2997/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2997/T5	I0/I2997/net13	I0/I2997/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2997/T2	BL5	net932	I0/I2997/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I114/T3	I0/I114/net049	net932	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I114/T4	vss	I0/I114/net13	I0/I114/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3070/T5	I0/I3070/net13	I0/I3070/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3070/T2	BL7	net934	I0/I3070/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3038/T3	I0/I3038/net049	net934	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3038/T4	vss	I0/I3038/net13	I0/I3038/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3038/T5	I0/I3038/net13	I0/I3038/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3038/T2	BL6	net934	I0/I3038/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3072/T5	I0/I3072/net13	I0/I3072/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3072/T2	BL7	net933	I0/I3072/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3040/T3	I0/I3040/net049	net933	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3040/T4	vss	I0/I3040/net13	I0/I3040/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3040/T5	I0/I3040/net13	I0/I3040/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3040/T2	BL6	net933	I0/I3040/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3061/T5	I0/I3061/net13	I0/I3061/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3061/T2	BL7	net932	I0/I3061/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3029/T3	I0/I3029/net049	net932	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3029/T4	vss	I0/I3029/net13	I0/I3029/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3029/T5	I0/I3029/net13	I0/I3029/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3029/T2	BL6	net932	I0/I3029/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2823/T3	I0/I2823/net049	net934	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2823/T4	vss	I0/I2823/net13	I0/I2823/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2823/T5	I0/I2823/net13	I0/I2823/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2823/T2	BL0	net934	I0/I2823/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3070/T3	I0/I3070/net049	net934	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3070/T4	vss	I0/I3070/net13	I0/I3070/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2824/T3	I0/I2824/net049	net933	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2824/T4	vss	I0/I2824/net13	I0/I2824/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2824/T5	I0/I2824/net13	I0/I2824/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2824/T2	BL0	net933	I0/I2824/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3072/T3	I0/I3072/net049	net933	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3072/T4	vss	I0/I3072/net13	I0/I3072/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2808/T3	I0/I2808/net049	net932	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2808/T4	vss	I0/I2808/net13	I0/I2808/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2808/T5	I0/I2808/net13	I0/I2808/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2808/T2	BL0	net932	I0/I2808/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3061/T3	I0/I3061/net049	net932	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3061/T4	vss	I0/I3061/net13	I0/I3061/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2897/T5	I0/I2897/net13	I0/I2897/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2897/T2	BL2	net934	I0/I2897/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2868/T3	I0/I2868/net049	net934	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2868/T4	vss	I0/I2868/net13	I0/I2868/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2868/T5	I0/I2868/net13	I0/I2868/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2868/T2	BL1	net934	I0/I2868/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2907/T5	I0/I2907/net13	I0/I2907/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2907/T2	BL2	net933	I0/I2907/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2874/T3	I0/I2874/net049	net933	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2874/T4	vss	I0/I2874/net13	I0/I2874/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2874/T5	I0/I2874/net13	I0/I2874/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2874/T2	BL1	net933	I0/I2874/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2917/T5	I0/I2917/net13	I0/I2917/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2917/T2	BL2	net932	I0/I2917/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2892/T3	I0/I2892/net049	net932	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2892/T4	vss	I0/I2892/net13	I0/I2892/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2892/T5	I0/I2892/net13	I0/I2892/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2892/T2	BL1	net932	I0/I2892/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2929/T3	I0/I2929/net049	net934	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2929/T4	vss	I0/I2929/net13	I0/I2929/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2929/T5	I0/I2929/net13	I0/I2929/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2929/T2	BL3	net934	I0/I2929/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2897/T3	I0/I2897/net049	net934	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2897/T4	vss	I0/I2897/net13	I0/I2897/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2945/T3	I0/I2945/net049	net933	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2945/T4	vss	I0/I2945/net13	I0/I2945/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2945/T5	I0/I2945/net13	I0/I2945/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2945/T2	BL3	net933	I0/I2945/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2907/T3	I0/I2907/net049	net933	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2907/T4	vss	I0/I2907/net13	I0/I2907/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2954/T3	I0/I2954/net049	net932	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2954/T4	vss	I0/I2954/net13	I0/I2954/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2954/T5	I0/I2954/net13	I0/I2954/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2954/T2	BL3	net932	I0/I2954/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2917/T3	I0/I2917/net049	net932	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2917/T4	vss	I0/I2917/net13	I0/I2917/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T431	net935	I1/net1944	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T441	net934	I1/net1972	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T448	net933	I1/net2000	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T434	I1/net864	I1/net1960	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T445	I1/net908	I1/net1984	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T454	I1/net944	I1/net2012	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T433	I1/net860	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T442	I1/net1972	I1/net908	I1/net900	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T443	I1/net900	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T449	I1/net2000	I1/net944	I1/net928	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T450	I1/net928	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T436	I1/net872	I1/a3bar	I1/net876	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T437	I1/net876	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T444	I1/net1984	I1/net880	I1/net912	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T446	I1/net912	I1/a3bar	I1/net916	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T447	I1/net916	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T451	I1/net2012	I1/net880	I1/net936	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T452	I1/net936	I1/a3	I1/net940	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T453	I1/net940	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T440	I1/net888	I1/a2	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T439	I1/net884	I1/a1bar	I1/net888	vss	nfet
+ L=0.12U	W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T438	I1/net880	I1/net1932	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T462	I1/net1932	I1/a0	I1/net884	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3171/T3	I0/I3171/net049	net931	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3171/T4	vss	I0/I3171/net13	I0/I3171/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3171/T5	I0/I3171/net13	I0/I3171/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3171/T2	BL10	net931	I0/I3171/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3139/T3	I0/I3139/net049	net931	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3139/T4	vss	I0/I3139/net13	I0/I3139/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3139/T5	I0/I3139/net13	I0/I3139/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3139/T2	BL9	net931	I0/I3139/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3107/T3	I0/I3107/net049	net931	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3107/T4	vss	I0/I3107/net13	I0/I3107/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3107/T5	I0/I3107/net13	I0/I3107/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3165/T3	I0/I3165/net049	net930	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3165/T4	vss	I0/I3165/net13	I0/I3165/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3165/T5	I0/I3165/net13	I0/I3165/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3165/T2	BL10	net930	I0/I3165/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3133/T3	I0/I3133/net049	net930	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3133/T4	vss	I0/I3133/net13	I0/I3133/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3133/T5	I0/I3133/net13	I0/I3133/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3133/T2	BL9	net930	I0/I3133/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3101/T3	I0/I3101/net049	net930	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3101/T4	vss	I0/I3101/net13	I0/I3101/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3101/T5	I0/I3101/net13	I0/I3101/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I100/T5	I0/I100/net13	I0/I100/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I100/T2	BL4	net931	I0/I100/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3203/T3	I0/I3203/net049	net931	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3203/T4	vss	I0/I3203/net13	I0/I3203/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3203/T5	I0/I3203/net13	I0/I3203/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3203/T2	BL11	net931	I0/I3203/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I106/T5	I0/I106/net13	I0/I106/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I106/T2	BL4	net930	I0/I106/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3197/T3	I0/I3197/net049	net930	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3197/T4	vss	I0/I3197/net13	I0/I3197/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3197/T5	I0/I3197/net13	I0/I3197/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3197/T2	BL11	net930	I0/I3197/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3011/T3	I0/I3011/net049	net931	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3011/T4	vss	I0/I3011/net13	I0/I3011/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3011/T5	I0/I3011/net13	I0/I3011/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3011/T2	BL5	net931	I0/I3011/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I100/T3	I0/I100/net049	net931	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I100/T4	vss	I0/I100/net13	I0/I100/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3005/T3	I0/I3005/net049	net930	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3005/T4	vss	I0/I3005/net13	I0/I3005/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3005/T5	I0/I3005/net13	I0/I3005/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3005/T2	BL5	net930	I0/I3005/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I106/T3	I0/I106/net049	net930	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I106/T4	vss	I0/I106/net13	I0/I106/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3075/T5	I0/I3075/net13	I0/I3075/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3075/T2	BL7	net931	I0/I3075/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3043/T3	I0/I3043/net049	net931	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3043/T4	vss	I0/I3043/net13	I0/I3043/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3043/T5	I0/I3043/net13	I0/I3043/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3043/T2	BL6	net931	I0/I3043/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3069/T5	I0/I3069/net13	I0/I3069/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3069/T2	BL7	net930	I0/I3069/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3037/T3	I0/I3037/net049	net930	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3037/T4	vss	I0/I3037/net13	I0/I3037/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3037/T5	I0/I3037/net13	I0/I3037/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3037/T2	BL6	net930	I0/I3037/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2819/T3	I0/I2819/net049	net931	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2819/T4	vss	I0/I2819/net13	I0/I2819/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2819/T5	I0/I2819/net13	I0/I2819/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2819/T2	BL0	net931	I0/I2819/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3075/T3	I0/I3075/net049	net931	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3075/T4	vss	I0/I3075/net13	I0/I3075/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2815/T3	I0/I2815/net049	net930	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2815/T4	vss	I0/I2815/net13	I0/I2815/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2815/T5	I0/I2815/net13	I0/I2815/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2815/T2	BL0	net930	I0/I2815/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3069/T3	I0/I3069/net049	net930	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3069/T4	vss	I0/I3069/net13	I0/I3069/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2924/T5	I0/I2924/net13	I0/I2924/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2924/T2	BL2	net931	I0/I2924/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2882/T3	I0/I2882/net049	net931	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2882/T4	vss	I0/I2882/net13	I0/I2882/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2882/T5	I0/I2882/net13	I0/I2882/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2882/T2	BL1	net931	I0/I2882/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2921/T5	I0/I2921/net13	I0/I2921/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2921/T2	BL2	net930	I0/I2921/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2873/T3	I0/I2873/net049	net930	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2873/T4	vss	I0/I2873/net13	I0/I2873/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2873/T5	I0/I2873/net13	I0/I2873/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2873/T2	BL1	net930	I0/I2873/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2955/T3	I0/I2955/net049	net931	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2955/T4	vss	I0/I2955/net13	I0/I2955/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2955/T5	I0/I2955/net13	I0/I2955/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2955/T2	BL3	net931	I0/I2955/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2924/T3	I0/I2924/net049	net931	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2924/T4	vss	I0/I2924/net13	I0/I2924/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2946/T3	I0/I2946/net049	net930	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2946/T4	vss	I0/I2946/net13	I0/I2946/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2946/T5	I0/I2946/net13	I0/I2946/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2946/T2	BL3	net930	I0/I2946/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2921/T3	I0/I2921/net049	net930	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2921/T4	vss	I0/I2921/net13	I0/I2921/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T461	net932	I1/net2044	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T526	net931	I1/net2096	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T455	I1/net948	I1/net2032	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T523	I1/net1076	I1/net1908	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T460	I1/net2044	I1/net948	I1/net964	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T459	I1/net964	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T525	I1/net2096	I1/net1076	I1/net1064	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T524	I1/net1064	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T519	I1/net1056	I1/net2136	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T458	I1/net2032	I1/net880	I1/net956	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T457	I1/net956	I1/a3	I1/net952	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T456	I1/net952	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T522	I1/net1908	I1/net1056	I1/net1104	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T521	I1/net1104	I1/a3bar	I1/net1060	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T520	I1/net1060	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3169/T3	I0/I3169/net049	net929	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3169/T4	vss	I0/I3169/net13	I0/I3169/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3169/T5	I0/I3169/net13	I0/I3169/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3169/T2	BL10	net929	I0/I3169/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3137/T3	I0/I3137/net049	net929	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3137/T4	vss	I0/I3137/net13	I0/I3137/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3137/T5	I0/I3137/net13	I0/I3137/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3137/T2	BL9	net929	I0/I3137/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3105/T3	I0/I3105/net049	net929	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3105/T4	vss	I0/I3105/net13	I0/I3105/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3105/T5	I0/I3105/net13	I0/I3105/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3181/T3	I0/I3181/net049	net928	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3181/T4	vss	I0/I3181/net13	I0/I3181/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3181/T5	I0/I3181/net13	I0/I3181/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3181/T2	BL10	net928	I0/I3181/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3149/T3	I0/I3149/net049	net928	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3149/T4	vss	I0/I3149/net13	I0/I3149/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3149/T5	I0/I3149/net13	I0/I3149/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3149/T2	BL9	net928	I0/I3149/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3117/T3	I0/I3117/net049	net928	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3117/T4	vss	I0/I3117/net13	I0/I3117/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3117/T5	I0/I3117/net13	I0/I3117/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I102/T5	I0/I102/net13	I0/I102/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I102/T2	BL4	net929	I0/I102/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3201/T3	I0/I3201/net049	net929	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3201/T4	vss	I0/I3201/net13	I0/I3201/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3201/T5	I0/I3201/net13	I0/I3201/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3201/T2	BL11	net929	I0/I3201/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I90/T5	I0/I90/net13	I0/I90/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I90/T2	BL4	net928	I0/I90/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3213/T3	I0/I3213/net049	net928	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3213/T4	vss	I0/I3213/net13	I0/I3213/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3213/T5	I0/I3213/net13	I0/I3213/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3213/T2	BL11	net928	I0/I3213/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3009/T3	I0/I3009/net049	net929	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3009/T4	vss	I0/I3009/net13	I0/I3009/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3009/T5	I0/I3009/net13	I0/I3009/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3009/T2	BL5	net929	I0/I3009/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I102/T3	I0/I102/net049	net929	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I102/T4	vss	I0/I102/net13	I0/I102/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3021/T3	I0/I3021/net049	net928	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3021/T4	vss	I0/I3021/net13	I0/I3021/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3021/T5	I0/I3021/net13	I0/I3021/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3021/T2	BL5	net928	I0/I3021/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I90/T3	I0/I90/net049	net928	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I90/T4	vss	I0/I90/net13	I0/I90/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3073/T5	I0/I3073/net13	I0/I3073/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3073/T2	BL7	net929	I0/I3073/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3041/T3	I0/I3041/net049	net929	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3041/T4	vss	I0/I3041/net13	I0/I3041/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3041/T5	I0/I3041/net13	I0/I3041/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3041/T2	BL6	net929	I0/I3041/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3085/T5	I0/I3085/net13	I0/I3085/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3085/T2	BL7	net928	I0/I3085/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3053/T3	I0/I3053/net049	net928	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3053/T4	vss	I0/I3053/net13	I0/I3053/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3053/T5	I0/I3053/net13	I0/I3053/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3053/T2	BL6	net928	I0/I3053/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2814/T3	I0/I2814/net049	net929	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2814/T4	vss	I0/I2814/net13	I0/I2814/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2814/T5	I0/I2814/net13	I0/I2814/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2814/T2	BL0	net929	I0/I2814/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3073/T3	I0/I3073/net049	net929	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3073/T4	vss	I0/I3073/net13	I0/I3073/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2818/T3	I0/I2818/net049	net928	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2818/T4	vss	I0/I2818/net13	I0/I2818/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2818/T5	I0/I2818/net13	I0/I2818/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2818/T2	BL0	net928	I0/I2818/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3085/T3	I0/I3085/net049	net928	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3085/T4	vss	I0/I3085/net13	I0/I3085/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2911/T5	I0/I2911/net13	I0/I2911/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2911/T2	BL2	net929	I0/I2911/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2876/T3	I0/I2876/net049	net929	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2876/T4	vss	I0/I2876/net13	I0/I2876/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2876/T5	I0/I2876/net13	I0/I2876/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2876/T2	BL1	net929	I0/I2876/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2898/T5	I0/I2898/net13	I0/I2898/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2898/T2	BL2	net928	I0/I2898/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2870/T3	I0/I2870/net049	net928	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2870/T4	vss	I0/I2870/net13	I0/I2870/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2870/T5	I0/I2870/net13	I0/I2870/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2870/T2	BL1	net928	I0/I2870/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2944/T3	I0/I2944/net049	net929	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2944/T4	vss	I0/I2944/net13	I0/I2944/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2944/T5	I0/I2944/net13	I0/I2944/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2944/T2	BL3	net929	I0/I2944/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2911/T3	I0/I2911/net049	net929	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2911/T4	vss	I0/I2911/net13	I0/I2911/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2930/T3	I0/I2930/net049	net928	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2930/T4	vss	I0/I2930/net13	I0/I2930/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2930/T5	I0/I2930/net13	I0/I2930/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2930/T2	BL3	net928	I0/I2930/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2898/T3	I0/I2898/net049	net928	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2898/T4	vss	I0/I2898/net13	I0/I2898/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T516	net930	I1/net2140	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T509	net929	I1/net1744	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T512	I1/net1116	I1/net1396	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T503	I1/net556	I1/net2120	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T515	I1/net2140	I1/net1116	I1/net1108	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T514	I1/net1108	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T508	I1/net1744	I1/net556	I1/net648	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T507	I1/net648	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T497	I1/net2152	I1/net560	I1/net1080	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T513	I1/net1396	I1/net1056	I1/net1124	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T511	I1/net1124	I1/a3bar	I1/net760	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T510	I1/net760	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T506	I1/net2120	I1/net1056	I1/net816	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T505	I1/net816	I1/a3	I1/net576	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T504	I1/net576	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T499	I1/net1892	I1/net1056	I1/net1068	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T99	vss	I1/net02030	I1/net02033	vss	nfet	L=0.12U
+ W=4.19U
+ AD=1.5503P	AS=1.5084P	PD=9.12U	PS=9.1U
+ wt=4.19e-06 wf=4.19e-06 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=5.748e-13 nrs=0.053076 nrd=0.053076 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T517	I1/net840	I1/a2bar	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T518	I1/net820	I1/a1	I1/net840	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T495	I1/net2136	I1/a0	I1/net820	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3135/T3	I0/I3135/net049	net927	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3135/T4	vss	I0/I3135/net13	I0/I3135/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3135/T5	I0/I3135/net13	I0/I3135/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3135/T2	BL9	net927	I0/I3135/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3103/T3	I0/I3103/net049	net927	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3103/T4	vss	I0/I3103/net13	I0/I3103/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3103/T5	I0/I3103/net13	I0/I3103/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3199/T4	vss	I0/I3199/net13	I0/I3199/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3199/T5	I0/I3199/net13	I0/I3199/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3199/T2	BL11	net927	I0/I3199/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3167/T3	I0/I3167/net049	net927	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3167/T4	vss	I0/I3167/net13	I0/I3167/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3167/T5	I0/I3167/net13	I0/I3167/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3167/T2	BL10	net927	I0/I3167/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3199/T3	I0/I3199/net049	net927	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3007/T4	vss	I0/I3007/net13	I0/I3007/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3007/T5	I0/I3007/net13	I0/I3007/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3007/T2	BL5	net927	I0/I3007/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I104/T3	I0/I104/net049	net927	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I104/T4	vss	I0/I104/net13	I0/I104/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I104/T5	I0/I104/net13	I0/I104/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I104/T2	BL4	net927	I0/I104/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3071/T2	BL7	net927	I0/I3071/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3039/T3	I0/I3039/net049	net927	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3039/T4	vss	I0/I3039/net13	I0/I3039/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3039/T5	I0/I3039/net13	I0/I3039/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3039/T2	BL6	net927	I0/I3039/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3007/T3	I0/I3007/net049	net927	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3146/T3	I0/I3146/net049	net926	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3146/T4	vss	I0/I3146/net13	I0/I3146/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3146/T5	I0/I3146/net13	I0/I3146/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3146/T2	BL9	net926	I0/I3146/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3114/T3	I0/I3114/net049	net926	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3114/T4	vss	I0/I3114/net13	I0/I3114/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3114/T5	I0/I3114/net13	I0/I3114/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3210/T4	vss	I0/I3210/net13	I0/I3210/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3210/T5	I0/I3210/net13	I0/I3210/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3210/T2	BL11	net926	I0/I3210/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3178/T3	I0/I3178/net049	net926	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3178/T4	vss	I0/I3178/net13	I0/I3178/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3178/T5	I0/I3178/net13	I0/I3178/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3178/T2	BL10	net926	I0/I3178/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3210/T3	I0/I3210/net049	net926	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3018/T4	vss	I0/I3018/net13	I0/I3018/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3018/T5	I0/I3018/net13	I0/I3018/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3018/T2	BL5	net926	I0/I3018/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I93/T3	I0/I93/net049	net926	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I93/T4	vss	I0/I93/net13	I0/I93/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I93/T5	I0/I93/net13	I0/I93/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I93/T2	BL4	net926	I0/I93/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3082/T2	BL7	net926	I0/I3082/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3050/T3	I0/I3050/net049	net926	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3050/T4	vss	I0/I3050/net13	I0/I3050/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3050/T5	I0/I3050/net13	I0/I3050/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3050/T2	BL6	net926	I0/I3050/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3018/T3	I0/I3018/net049	net926	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3145/T3	I0/I3145/net049	net925	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3145/T4	vss	I0/I3145/net13	I0/I3145/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3145/T5	I0/I3145/net13	I0/I3145/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3145/T2	BL9	net925	I0/I3145/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3113/T3	I0/I3113/net049	net925	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3113/T4	vss	I0/I3113/net13	I0/I3113/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3113/T5	I0/I3113/net13	I0/I3113/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3209/T4	vss	I0/I3209/net13	I0/I3209/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3209/T5	I0/I3209/net13	I0/I3209/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3209/T2	BL11	net925	I0/I3209/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3177/T3	I0/I3177/net049	net925	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3177/T4	vss	I0/I3177/net13	I0/I3177/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3177/T5	I0/I3177/net13	I0/I3177/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3177/T2	BL10	net925	I0/I3177/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3209/T3	I0/I3209/net049	net925	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3017/T4	vss	I0/I3017/net13	I0/I3017/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3017/T5	I0/I3017/net13	I0/I3017/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3017/T2	BL5	net925	I0/I3017/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I94/T3	I0/I94/net049	net925	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I94/T4	vss	I0/I94/net13	I0/I94/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I94/T5	I0/I94/net13	I0/I94/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I94/T2	BL4	net925	I0/I94/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3081/T2	BL7	net925	I0/I3081/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3049/T3	I0/I3049/net049	net925	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3049/T4	vss	I0/I3049/net13	I0/I3049/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3049/T5	I0/I3049/net13	I0/I3049/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3049/T2	BL6	net925	I0/I3049/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3017/T3	I0/I3017/net049	net925	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3122/T3	I0/I3122/net049	net924	BL9bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3122/T4	vss	I0/I3122/net13	I0/I3122/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3122/T5	I0/I3122/net13	I0/I3122/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3122/T2	BL9	net924	I0/I3122/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3090/T3	I0/I3090/net049	net924	BL8bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3090/T4	vss	I0/I3090/net13	I0/I3090/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3090/T5	I0/I3090/net13	I0/I3090/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3186/T4	vss	I0/I3186/net13	I0/I3186/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3186/T5	I0/I3186/net13	I0/I3186/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3186/T2	BL11	net924	I0/I3186/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3154/T3	I0/I3154/net049	net924	BL10bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3154/T4	vss	I0/I3154/net13	I0/I3154/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3154/T5	I0/I3154/net13	I0/I3154/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3154/T2	BL10	net924	I0/I3154/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3186/T3	I0/I3186/net049	net924	BL11bar	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2994/T4	vss	I0/I2994/net13	I0/I2994/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2994/T5	I0/I2994/net13	I0/I2994/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2994/T2	BL5	net924	I0/I2994/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I117/T3	I0/I117/net049	net924	BL4bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I117/T4	vss	I0/I117/net13	I0/I117/net049	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I117/T5	I0/I117/net13	I0/I117/net049	vss	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I117/T2	BL4	net924	I0/I117/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3058/T2	BL7	net924	I0/I3058/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3026/T3	I0/I3026/net049	net924	BL6bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3026/T4	vss	I0/I3026/net13	I0/I3026/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3026/T5	I0/I3026/net13	I0/I3026/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3026/T2	BL6	net924	I0/I3026/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2994/T3	I0/I2994/net049	net924	BL5bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI52/T1	net741	y4	BL11bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI53/T1	BL11	y4	net740	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI54/T1	net741	y3	BL10bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI55/T1	BL10	y3	net740	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI56/T1	net741	y2	BL9bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI57/T1	BL9	y2	net740	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI58/T1	net741	y1	BL8bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T4	vss	vdd	I22/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T8	vss	I22/net20	I22/net8	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T7	data0	I22/net8	vss	vss	nfet	L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T11	I23/net23	data0	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T16	I23/net15	net680	net220	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.32P	PD=1.36U	PS=2.64U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T17	vss	I23/net23	I23/net15	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T19	I23/net7	net220	vss	vss	nfet	L=0.12U
+ W=1U
+ AD=0.18P	AS=0.18P	PD=1.36U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T18	net208	net680	I23/net7	vss	nfet	L=0.12U
+ W=1U
+ AD=0.32P	AS=0.18P	PD=2.64U	PS=1.36U
+ wt=1e-06 wf=1e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.230366 nrd=0.230366 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T2	I2/net23	net262	I2/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T3	I2/net20	net256	I2/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T4	vss	vdd	I2/net23	vss	nfet	L=0.12U	W=5U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.12e-14 panw8=2.4e-14 panw7=1.2e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI45/T1	BL7	y4	net262	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI46/T1	net256	y3	BL6bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI47/T1	BL6	y3	net262	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI48/T1	net256	y2	BL5bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI49/T1	BL5	y2	net262	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI50/T1	net256	y1	BL4bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T2	I22/net23	net220	I22/net24	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI51/T1	BL4	y1	net262	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T3	I22/net20	net208	I22/net23	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.16e-14 panw7=1.2e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T65	y4bar	I116/net0113	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.796e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T67	I116/net0101	I116/net0105	vss	vss	nfet	L=0.12U
+ W=1.18U
+ AD=0.3776P	AS=0.3776P	PD=3U	PS=3U
+ wt=1.18e-06 wf=1.18e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.59e-13 panw8=5.94e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.193833 nrd=0.193833 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI30/T22	vss	I30/net41	net680	vss	nfet	L=0.12U
+ W=4.5U
+ AD=1.44P	AS=1.44P	PD=9.64U	PS=9.64U
+ wt=4.5e-06 wf=4.5e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.368e-13 panw7=4.032e-13 nrs=0.0493827 nrd=0.0493827 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI30/T21	I30/net41	I30/net17	vss	vss	nfet	L=0.12U
+ W=1.22U
+ AD=0.3904P	AS=0.3904P	PD=3.08U	PS=3.08U
+ wt=1.22e-06 wf=1.22e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.704e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-14 nrs=0.187234 nrd=0.187234 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T496	net928	I1/net2152	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.02e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2869/T5	I0/I2869/net13	I0/I2869/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2869/T2	BL1	net927	I0/I2869/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2822/T3	I0/I2822/net049	net927	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2822/T4	vss	I0/I2822/net13	I0/I2822/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2822/T5	I0/I2822/net13	I0/I2822/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2822/T2	BL0	net927	I0/I2822/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3071/T3	I0/I3071/net049	net927	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3071/T4	vss	I0/I3071/net13	I0/I3071/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3071/T5	I0/I3071/net13	I0/I3071/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2869/T4	vss	I0/I2869/net13	I0/I2869/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2931/T3	I0/I2931/net049	net927	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2931/T4	vss	I0/I2931/net13	I0/I2931/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2931/T5	I0/I2931/net13	I0/I2931/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2931/T2	BL3	net927	I0/I2931/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2899/T3	I0/I2899/net049	net927	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2899/T4	vss	I0/I2899/net13	I0/I2899/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2899/T5	I0/I2899/net13	I0/I2899/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2899/T2	BL2	net927	I0/I2899/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2869/T3	I0/I2869/net049	net927	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2878/T5	I0/I2878/net13	I0/I2878/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2878/T2	BL1	net926	I0/I2878/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2817/T3	I0/I2817/net049	net926	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2817/T4	vss	I0/I2817/net13	I0/I2817/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2817/T5	I0/I2817/net13	I0/I2817/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2817/T2	BL0	net926	I0/I2817/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3082/T3	I0/I3082/net049	net926	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3082/T4	vss	I0/I3082/net13	I0/I3082/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3082/T5	I0/I3082/net13	I0/I3082/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2878/T4	vss	I0/I2878/net13	I0/I2878/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2927/T3	I0/I2927/net049	net926	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2927/T4	vss	I0/I2927/net13	I0/I2927/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2927/T5	I0/I2927/net13	I0/I2927/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2927/T2	BL3	net926	I0/I2927/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2900/T3	I0/I2900/net049	net926	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2900/T4	vss	I0/I2900/net13	I0/I2900/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2900/T5	I0/I2900/net13	I0/I2900/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2900/T2	BL2	net926	I0/I2900/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2878/T3	I0/I2878/net049	net926	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T559	net927	I1/net2060	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.95e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2806/T3	I0/I2806/net049	net925	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2806/T4	vss	I0/I2806/net13	I0/I2806/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2806/T5	I0/I2806/net13	I0/I2806/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2806/T2	BL0	net925	I0/I2806/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3081/T3	I0/I3081/net049	net925	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3081/T4	vss	I0/I3081/net13	I0/I3081/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3081/T5	I0/I3081/net13	I0/I3081/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2904/T4	vss	I0/I2904/net13	I0/I2904/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2904/T5	I0/I2904/net13	I0/I2904/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2904/T2	BL2	net925	I0/I2904/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2884/T3	I0/I2884/net049	net925	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2884/T4	vss	I0/I2884/net13	I0/I2884/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2884/T5	I0/I2884/net13	I0/I2884/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2884/T2	BL1	net925	I0/I2884/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2904/T3	I0/I2904/net049	net925	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T569	net926	I1/net2212	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I2939/T3	I0/I2939/net049	net925	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2939/T4	vss	I0/I2939/net13	I0/I2939/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2939/T5	I0/I2939/net13	I0/I2939/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2939/T2	BL3	net925	I0/I2939/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2863/T5	I0/I2863/net13	I0/I2863/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2863/T2	BL1	net924	I0/I2863/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2807/T3	I0/I2807/net049	net924	BL0bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2807/T4	vss	I0/I2807/net13	I0/I2807/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2807/T5	I0/I2807/net13	I0/I2807/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2807/T2	BL0	net924	I0/I2807/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3058/T3	I0/I3058/net049	net924	BL7bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3058/T4	vss	I0/I3058/net13	I0/I3058/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3058/T5	I0/I3058/net13	I0/I3058/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2863/T4	vss	I0/I2863/net13	I0/I2863/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2937/T3	I0/I2937/net049	net924	BL3bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2937/T4	vss	I0/I2937/net13	I0/I2937/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2937/T5	I0/I2937/net13	I0/I2937/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2937/T2	BL3	net924	I0/I2937/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2925/T3	I0/I2925/net049	net924	BL2bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2925/T4	vss	I0/I2925/net13	I0/I2925/net049	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2925/T5	I0/I2925/net13	I0/I2925/net049	vss	vss	nfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0504P	PD=0.64U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2925/T2	BL2	net924	I0/I2925/net13	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2863/T3	I0/I2863/net049	net924	BL1bar	vss	nfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T576	net925	I1/net2068	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.23e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI37/T1	net208	y1	BL0bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T69	I116/net0229	I116/net0373	I116/net0282	vss	nfet
+ L=0.12U	W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26U	PS=1.17U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.452e-13 panw8=2.4e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T80	I116/net0282	I116/net56	vss	vss	nfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17U	PS=2.26U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=9.72e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI36/T1	BL0	y1	net220	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T66	vss	I116/net0229	I116/net0105	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI44/T1	net256	y4	BL7bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T68	y4	I116/net0101	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=1.003e-13 panw7=7.85e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI41/T1	net208	y3	BL2bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T9	I116/net56	I116/net60	vss	vss	nfet	L=0.12U
+ W=0.6U
+ AD=0.192P	AS=0.192P	PD=1.84U	PS=1.84U
+ wt=6e-07 wf=6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI40/T1	BL2	y3	net220	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T64	vss	I116/net0229	I116/net0113	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=7.32e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI39/T1	net208	y2	BL1bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI38/T1	BL1	y2	net220	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T54	vss	I116/net0281	I116/net0125	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=7.68e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T589	net924	I1/net2224	vss	vss	nfet	L=0.12U
+ W=3.62U
+ AD=1.3032P	AS=1.3394P	PD=7.96U	PS=7.98U
+ wt=3.62e-06 wf=3.62e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=1.332e-13 nrs=0.0615385 nrd=0.0615385 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T52	vss	I116/net0281	I116/net0133	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T50	y3	I116/net0137	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=1.003e-13 panw7=7.85e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.236e-13 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T8	I116/net60	addr6	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T49	I116/net0281	I116/net120	I116/net0286	vss	nfet
+ L=0.12U	W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26U	PS=1.17U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.332e-13 panw8=2.4e-14 panw7=1.2e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T79	I116/net0286	I116/net0373	vss	vss	nfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17U	PS=2.26U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=9.72e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI43/T1	net208	y4	BL3bar	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI42/T1	BL3	y4	net220	vss	nfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=8.4e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T53	y3bar	I116/net0125	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.796e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T502	I1/net560	I1/net1892	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T562	I1/net1008	I1/net2256	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T573	I1/net1152	I1/net2216	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T582	I1/net1000	I1/net2192	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T498	I1/net1080	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T560	I1/net2060	I1/net1008	I1/net1012	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T561	I1/net1012	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T570	I1/net2212	I1/net1152	I1/net1156	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T571	I1/net1156	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T577	I1/net2068	I1/net1000	I1/net1020	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T578	I1/net1020	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T583	I1/net1132	I1/net2236	vss	vss	nfet	L=0.12U
+ W=0.56U
+ AD=0.2016P	AS=0.2072P	PD=1.84U	PS=1.86U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=9.6e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T588	I1/net2224	I1/net1132	I1/net848	vss	nfet
+ L=0.12U	W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T587	I1/net848	I1/addr_en_b	vss	vss	nfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.16e-14 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T11	I116/net0373	I116/net52	vss	vss	nfet	L=0.12U
+ W=0.6U
+ AD=0.192P	AS=0.192P	PD=1.84U	PS=1.84U
+ wt=6e-07 wf=6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=6.8e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T2	I116/net120	addr6	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T25	vss	I116/net96	I116/net24	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=7.68e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T7	I116/net116	addr5	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T12	I116/net96	I116/net116	I116/net0342	vss	nfet
+ L=0.12U	W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26U	PS=1.17U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.332e-13 panw8=2.4e-14 panw7=1.2e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T77	I116/net0342	I116/net120	vss	vss	nfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17U	PS=2.26U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=9.72e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T22	vss	I116/net96	I116/net32	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T20	y1	I116/net36	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=1.003e-13 panw7=7.85e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.236e-13 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T23	y1bar	I116/net24	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.796e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T21	I116/net36	I116/net32	vss	vss	nfet	L=0.12U
+ W=1.18U
+ AD=0.3776P	AS=0.3776P	PD=3U	PS=3U
+ wt=1.18e-06 wf=1.18e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.638e-13 panw8=5.94e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.193833 nrd=0.193833 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T51	I116/net0137	I116/net0133	vss	vss	nfet	L=0.12U
+ W=1.18U
+ AD=0.3776P	AS=0.3776P	PD=3U	PS=3U
+ wt=1.18e-06 wf=1.18e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw10=9.44e-14 nrs=0.193833 nrd=0.193833 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T36	vss	I116/net0309	I116/net0157	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=7.68e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T500	I1/net1068	I1/a3	I1/net1072	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T501	I1/net1072	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T563	I1/net2256	I1/net612	I1/net996	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T564	I1/net996	I1/a3bar	I1/net1128	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T565	I1/net1128	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T572	I1/net2216	I1/net612	I1/net1036	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T574	I1/net1036	I1/a3bar	I1/net1032	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T575	I1/net1032	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T579	I1/net2192	I1/net612	I1/net1004	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T580	I1/net1004	I1/a3	I1/net1136	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T568	I1/net1048	I1/a2	vss	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0814P	AS=0.1408P	PD=0.81U	PS=1.52U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T567	I1/net592	I1/a1	I1/net1048	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.0792P	AS=0.0814P	PD=0.8U	PS=0.81U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T566	I1/net612	I1/net2184	vss	vss	nfet	L=0.12U
+ W=0.43U
+ AD=0.1548P	AS=0.1591P	PD=1.58U	PS=1.6U
+ wt=4.3e-07 wf=4.3e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=1.56e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.571429 nrd=0.571429 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T590	I1/net2184	I1/a0	I1/net592	vss	nfet	L=0.12U
+ W=0.44U
+ AD=0.1408P	AS=0.0792P	PD=1.52U	PS=0.8U
+ wt=4.4e-07 wf=4.4e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.556962 nrd=0.556962 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T38	vss	I116/net0309	I116/net0149	vss	nfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T40	y2	I116/net0145	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=1.003e-13 panw7=7.85e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.236e-13 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T10	I116/net52	addr5	vss	vss	nfet	L=0.12U
+ W=0.33U
+ AD=0.1056P	AS=0.1056P	PD=1.3U	PS=1.3U
+ wt=3.3e-07 wf=3.3e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.77193 nrd=0.77193 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T581	I1/net1136	I1/a4bar	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T586	I1/net2236	I1/net612	I1/net980	vss	nfet
+ L=0.12U	W=0.57U
+ AD=0.1824P	AS=0.1026P	PD=1.78U	PS=0.93U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T585	I1/net980	I1/a3	I1/net984	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.1026P	AS=0.10545P	PD=0.93U	PS=0.94U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T584	I1/net984	I1/a4	vss	vss	nfet	L=0.12U
+ W=0.57U
+ AD=0.10545P	AS=0.1824P	PD=0.94U	PS=1.78U
+ wt=5.7e-07 wf=5.7e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.52e-14 panw8=2.4e-14 panw7=1.92e-14 nrs=0.419048 nrd=0.419048 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T41	I116/net0309	I116/net116	I116/net0326	vss	nfet
+ L=0.12U	W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26U	PS=1.17U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.332e-13 panw8=2.4e-14 panw7=1.2e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T78	I116/net0326	I116/net56	vss	vss	nfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17U	PS=2.26U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=9.72e-14 panw10=2.52e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T37	y2bar	I116/net0157	vss	vss	nfet	L=0.12U
+ W=2.13U
+ AD=0.6816P	AS=0.6816P	PD=4.9U	PS=4.9U
+ wt=2.13e-06 wf=2.13e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.796e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.105516 nrd=0.105516 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T100	vss	I1/net02033	I1/addr_en_b	vss	nfet	L=0.12U
+ W=14.8U
+ AD=5.476P	AS=5.328P	PD=30.34U	PS=30.32U
+ wt=1.48e-05 wf=1.48e-05 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0149102 nrd=0.0149102 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T39	I116/net0145	I116/net0149	vss	vss	nfet	L=0.12U
+ W=1.18U
+ AD=0.3776P	AS=0.3776P	PD=3U	PS=3U
+ wt=1.18e-06 wf=1.18e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.506e-13 panw8=5.82e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=9.6e-15 nrs=0.193833 nrd=0.193833 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI156/T1	vdd	clkout	BL37bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4156/T0	vdd	I0/I4156/net13	I0/I4156/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI156/T2	BL37	clkout	BL37bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI156/T0	BL37	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4156/T1	I0/I4156/net13	I0/I4156/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI155/T1	vdd	clkout	BL36bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.464e-13 panw10=2.256e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4060/T0	vdd	I0/I4060/net13	I0/I4060/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.68e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.68e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI155/T2	BL36	clkout	BL36bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=7.2e-14 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI155/T0	BL36	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw8=2.4e-13 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4060/T1	I0/I4060/net13	I0/I4060/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI158/T0	BL39	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4220/T1	I0/I4220/net13	I0/I4220/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI157/T1	vdd	clkout	BL38bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4188/T0	vdd	I0/I4188/net13	I0/I4188/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI157/T2	BL38	clkout	BL38bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI157/T0	BL38	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4188/T1	I0/I4188/net13	I0/I4188/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI158/T2	BL39	clkout	BL39bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI151/T1	vdd	clkout	BL32bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3932/T0	vdd	I0/I3932/net13	I0/I3932/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI151/T2	BL32	clkout	BL32bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI151/T0	BL32	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3932/T1	I0/I3932/net13	I0/I3932/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI158/T1	vdd	clkout	BL39bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4220/T0	vdd	I0/I4220/net13	I0/I4220/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI153/T1	vdd	clkout	BL34bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3996/T0	vdd	I0/I3996/net13	I0/I3996/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI153/T2	BL34	clkout	BL34bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI153/T0	BL34	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3996/T1	I0/I3996/net13	I0/I3996/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI152/T1	vdd	clkout	BL33bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3964/T0	vdd	I0/I3964/net13	I0/I3964/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI152/T2	BL33	clkout	BL33bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI152/T0	BL33	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3964/T1	I0/I3964/net13	I0/I3964/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4148/T0	vdd	I0/I4148/net13	I0/I4148/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4147/T0	vdd	I0/I4147/net13	I0/I4147/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4148/T1	I0/I4148/net13	I0/I4148/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4147/T1	I0/I4147/net13	I0/I4147/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4052/T0	vdd	I0/I4052/net13	I0/I4052/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.68e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.68e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4051/T0	vdd	I0/I4051/net13	I0/I4051/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.68e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.68e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4052/T1	I0/I4052/net13	I0/I4052/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4051/T1	I0/I4051/net13	I0/I4051/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4212/T1	I0/I4212/net13	I0/I4212/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4211/T1	I0/I4211/net13	I0/I4211/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4180/T0	vdd	I0/I4180/net13	I0/I4180/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4179/T0	vdd	I0/I4179/net13	I0/I4179/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4180/T1	I0/I4180/net13	I0/I4180/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4179/T1	I0/I4179/net13	I0/I4179/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3924/T0	vdd	I0/I3924/net13	I0/I3924/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3923/T0	vdd	I0/I3923/net13	I0/I3923/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3924/T1	I0/I3924/net13	I0/I3924/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3923/T1	I0/I3923/net13	I0/I3923/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4212/T0	vdd	I0/I4212/net13	I0/I4212/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4211/T0	vdd	I0/I4211/net13	I0/I4211/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3988/T0	vdd	I0/I3988/net13	I0/I3988/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3987/T0	vdd	I0/I3987/net13	I0/I3987/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3988/T1	I0/I3988/net13	I0/I3988/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3987/T1	I0/I3987/net13	I0/I3987/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3956/T0	vdd	I0/I3956/net13	I0/I3956/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3955/T0	vdd	I0/I3955/net13	I0/I3955/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3956/T1	I0/I3956/net13	I0/I3956/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3955/T1	I0/I3955/net13	I0/I3955/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4076/T0	vdd	I0/I4076/net13	I0/I4076/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.68e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.68e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4057/T0	vdd	I0/I4057/net13	I0/I4057/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.68e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.68e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4072/T0	vdd	I0/I4072/net13	I0/I4072/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.12e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.24e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4070/T0	vdd	I0/I4070/net13	I0/I4070/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.12e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.24e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4076/T1	I0/I4076/net13	I0/I4076/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4057/T1	I0/I4057/net13	I0/I4057/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4072/T1	I0/I4072/net13	I0/I4072/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4070/T1	I0/I4070/net13	I0/I4070/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4172/T0	vdd	I0/I4172/net13	I0/I4172/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4153/T0	vdd	I0/I4153/net13	I0/I4153/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4168/T0	vdd	I0/I4168/net13	I0/I4168/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4166/T0	vdd	I0/I4166/net13	I0/I4166/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4172/T1	I0/I4172/net13	I0/I4172/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4153/T1	I0/I4153/net13	I0/I4153/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4168/T1	I0/I4168/net13	I0/I4168/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4166/T1	I0/I4166/net13	I0/I4166/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4204/T0	vdd	I0/I4204/net13	I0/I4204/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4185/T0	vdd	I0/I4185/net13	I0/I4185/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4200/T0	vdd	I0/I4200/net13	I0/I4200/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4198/T0	vdd	I0/I4198/net13	I0/I4198/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4204/T1	I0/I4204/net13	I0/I4204/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4185/T1	I0/I4185/net13	I0/I4185/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4200/T1	I0/I4200/net13	I0/I4200/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4198/T1	I0/I4198/net13	I0/I4198/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4236/T1	I0/I4236/net13	I0/I4236/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4217/T1	I0/I4217/net13	I0/I4217/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4232/T1	I0/I4232/net13	I0/I4232/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4230/T1	I0/I4230/net13	I0/I4230/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4236/T0	vdd	I0/I4236/net13	I0/I4236/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4217/T0	vdd	I0/I4217/net13	I0/I4217/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4232/T0	vdd	I0/I4232/net13	I0/I4232/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4230/T0	vdd	I0/I4230/net13	I0/I4230/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3948/T0	vdd	I0/I3948/net13	I0/I3948/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3929/T0	vdd	I0/I3929/net13	I0/I3929/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3944/T0	vdd	I0/I3944/net13	I0/I3944/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3942/T0	vdd	I0/I3942/net13	I0/I3942/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3948/T1	I0/I3948/net13	I0/I3948/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3929/T1	I0/I3929/net13	I0/I3929/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3944/T1	I0/I3944/net13	I0/I3944/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3942/T1	I0/I3942/net13	I0/I3942/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3980/T0	vdd	I0/I3980/net13	I0/I3980/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3961/T0	vdd	I0/I3961/net13	I0/I3961/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3976/T0	vdd	I0/I3976/net13	I0/I3976/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3974/T0	vdd	I0/I3974/net13	I0/I3974/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3980/T1	I0/I3980/net13	I0/I3980/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3961/T1	I0/I3961/net13	I0/I3961/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3976/T1	I0/I3976/net13	I0/I3976/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3974/T1	I0/I3974/net13	I0/I3974/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4012/T0	vdd	I0/I4012/net13	I0/I4012/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3993/T0	vdd	I0/I3993/net13	I0/I3993/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4008/T0	vdd	I0/I4008/net13	I0/I4008/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4006/T0	vdd	I0/I4006/net13	I0/I4006/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4012/T1	I0/I4012/net13	I0/I4012/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3993/T1	I0/I3993/net13	I0/I3993/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4008/T1	I0/I4008/net13	I0/I4008/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4006/T1	I0/I4006/net13	I0/I4006/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4066/T1	I0/I4066/net13	I0/I4066/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4058/T1	I0/I4058/net13	I0/I4058/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4059/T1	I0/I4059/net13	I0/I4059/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4049/T1	I0/I4049/net13	I0/I4049/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4075/T1	I0/I4075/net13	I0/I4075/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4069/T1	I0/I4069/net13	I0/I4069/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4055/T1	I0/I4055/net13	I0/I4055/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4048/T1	I0/I4048/net13	I0/I4048/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4071/T1	I0/I4071/net13	I0/I4071/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4068/T1	I0/I4068/net13	I0/I4068/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4066/T0	vdd	I0/I4066/net13	I0/I4066/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4058/T0	vdd	I0/I4058/net13	I0/I4058/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4059/T0	vdd	I0/I4059/net13	I0/I4059/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4049/T0	vdd	I0/I4049/net13	I0/I4049/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4075/T0	vdd	I0/I4075/net13	I0/I4075/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4069/T0	vdd	I0/I4069/net13	I0/I4069/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4055/T0	vdd	I0/I4055/net13	I0/I4055/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4048/T0	vdd	I0/I4048/net13	I0/I4048/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4071/T0	vdd	I0/I4071/net13	I0/I4071/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4068/T0	vdd	I0/I4068/net13	I0/I4068/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4162/T1	I0/I4162/net13	I0/I4162/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4154/T1	I0/I4154/net13	I0/I4154/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4155/T1	I0/I4155/net13	I0/I4155/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4145/T1	I0/I4145/net13	I0/I4145/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4171/T1	I0/I4171/net13	I0/I4171/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4165/T1	I0/I4165/net13	I0/I4165/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4151/T1	I0/I4151/net13	I0/I4151/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4144/T1	I0/I4144/net13	I0/I4144/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4167/T1	I0/I4167/net13	I0/I4167/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4164/T1	I0/I4164/net13	I0/I4164/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4162/T0	vdd	I0/I4162/net13	I0/I4162/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4154/T0	vdd	I0/I4154/net13	I0/I4154/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4155/T0	vdd	I0/I4155/net13	I0/I4155/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4145/T0	vdd	I0/I4145/net13	I0/I4145/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4171/T0	vdd	I0/I4171/net13	I0/I4171/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4165/T0	vdd	I0/I4165/net13	I0/I4165/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4151/T0	vdd	I0/I4151/net13	I0/I4151/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4144/T0	vdd	I0/I4144/net13	I0/I4144/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4167/T0	vdd	I0/I4167/net13	I0/I4167/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4164/T0	vdd	I0/I4164/net13	I0/I4164/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4194/T1	I0/I4194/net13	I0/I4194/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4186/T1	I0/I4186/net13	I0/I4186/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4187/T1	I0/I4187/net13	I0/I4187/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4177/T1	I0/I4177/net13	I0/I4177/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4203/T1	I0/I4203/net13	I0/I4203/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4197/T1	I0/I4197/net13	I0/I4197/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4183/T1	I0/I4183/net13	I0/I4183/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4176/T1	I0/I4176/net13	I0/I4176/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4199/T1	I0/I4199/net13	I0/I4199/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4196/T1	I0/I4196/net13	I0/I4196/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4194/T0	vdd	I0/I4194/net13	I0/I4194/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4186/T0	vdd	I0/I4186/net13	I0/I4186/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4187/T0	vdd	I0/I4187/net13	I0/I4187/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4177/T0	vdd	I0/I4177/net13	I0/I4177/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4203/T0	vdd	I0/I4203/net13	I0/I4203/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4197/T0	vdd	I0/I4197/net13	I0/I4197/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4183/T0	vdd	I0/I4183/net13	I0/I4183/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4176/T0	vdd	I0/I4176/net13	I0/I4176/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4199/T0	vdd	I0/I4199/net13	I0/I4199/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4196/T0	vdd	I0/I4196/net13	I0/I4196/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4226/T1	I0/I4226/net13	I0/I4226/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4218/T1	I0/I4218/net13	I0/I4218/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4219/T1	I0/I4219/net13	I0/I4219/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4209/T1	I0/I4209/net13	I0/I4209/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4235/T1	I0/I4235/net13	I0/I4235/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4229/T1	I0/I4229/net13	I0/I4229/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4215/T1	I0/I4215/net13	I0/I4215/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4208/T1	I0/I4208/net13	I0/I4208/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4231/T1	I0/I4231/net13	I0/I4231/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4228/T1	I0/I4228/net13	I0/I4228/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4226/T0	vdd	I0/I4226/net13	I0/I4226/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4218/T0	vdd	I0/I4218/net13	I0/I4218/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4219/T0	vdd	I0/I4219/net13	I0/I4219/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4209/T0	vdd	I0/I4209/net13	I0/I4209/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4235/T0	vdd	I0/I4235/net13	I0/I4235/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4229/T0	vdd	I0/I4229/net13	I0/I4229/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4215/T0	vdd	I0/I4215/net13	I0/I4215/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4208/T0	vdd	I0/I4208/net13	I0/I4208/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4231/T0	vdd	I0/I4231/net13	I0/I4231/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4228/T0	vdd	I0/I4228/net13	I0/I4228/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3938/T1	I0/I3938/net13	I0/I3938/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3930/T1	I0/I3930/net13	I0/I3930/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3931/T1	I0/I3931/net13	I0/I3931/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3921/T1	I0/I3921/net13	I0/I3921/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3947/T1	I0/I3947/net13	I0/I3947/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3941/T1	I0/I3941/net13	I0/I3941/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3927/T1	I0/I3927/net13	I0/I3927/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3920/T1	I0/I3920/net13	I0/I3920/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3943/T1	I0/I3943/net13	I0/I3943/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3940/T1	I0/I3940/net13	I0/I3940/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3938/T0	vdd	I0/I3938/net13	I0/I3938/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3930/T0	vdd	I0/I3930/net13	I0/I3930/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3931/T0	vdd	I0/I3931/net13	I0/I3931/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3921/T0	vdd	I0/I3921/net13	I0/I3921/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3947/T0	vdd	I0/I3947/net13	I0/I3947/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3941/T0	vdd	I0/I3941/net13	I0/I3941/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3927/T0	vdd	I0/I3927/net13	I0/I3927/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3920/T0	vdd	I0/I3920/net13	I0/I3920/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3943/T0	vdd	I0/I3943/net13	I0/I3943/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3940/T0	vdd	I0/I3940/net13	I0/I3940/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3970/T1	I0/I3970/net13	I0/I3970/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3962/T1	I0/I3962/net13	I0/I3962/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3963/T1	I0/I3963/net13	I0/I3963/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3953/T1	I0/I3953/net13	I0/I3953/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3979/T1	I0/I3979/net13	I0/I3979/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3973/T1	I0/I3973/net13	I0/I3973/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3959/T1	I0/I3959/net13	I0/I3959/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3952/T1	I0/I3952/net13	I0/I3952/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3975/T1	I0/I3975/net13	I0/I3975/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3972/T1	I0/I3972/net13	I0/I3972/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3970/T0	vdd	I0/I3970/net13	I0/I3970/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3962/T0	vdd	I0/I3962/net13	I0/I3962/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3963/T0	vdd	I0/I3963/net13	I0/I3963/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3953/T0	vdd	I0/I3953/net13	I0/I3953/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3979/T0	vdd	I0/I3979/net13	I0/I3979/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3973/T0	vdd	I0/I3973/net13	I0/I3973/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3959/T0	vdd	I0/I3959/net13	I0/I3959/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3952/T0	vdd	I0/I3952/net13	I0/I3952/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3975/T0	vdd	I0/I3975/net13	I0/I3975/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3972/T0	vdd	I0/I3972/net13	I0/I3972/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4002/T1	I0/I4002/net13	I0/I4002/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3994/T1	I0/I3994/net13	I0/I3994/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3995/T1	I0/I3995/net13	I0/I3995/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3985/T1	I0/I3985/net13	I0/I3985/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4011/T1	I0/I4011/net13	I0/I4011/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4005/T1	I0/I4005/net13	I0/I4005/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3991/T1	I0/I3991/net13	I0/I3991/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3984/T1	I0/I3984/net13	I0/I3984/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4007/T1	I0/I4007/net13	I0/I4007/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4004/T1	I0/I4004/net13	I0/I4004/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4002/T0	vdd	I0/I4002/net13	I0/I4002/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3994/T0	vdd	I0/I3994/net13	I0/I3994/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3995/T0	vdd	I0/I3995/net13	I0/I3995/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3985/T0	vdd	I0/I3985/net13	I0/I3985/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4011/T0	vdd	I0/I4011/net13	I0/I4011/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4005/T0	vdd	I0/I4005/net13	I0/I4005/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3991/T0	vdd	I0/I3991/net13	I0/I3991/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3984/T0	vdd	I0/I3984/net13	I0/I3984/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4007/T0	vdd	I0/I4007/net13	I0/I4007/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4004/T0	vdd	I0/I4004/net13	I0/I4004/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4046/T1	I0/I4046/net13	I0/I4046/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4047/T1	I0/I4047/net13	I0/I4047/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4054/T1	I0/I4054/net13	I0/I4054/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4056/T1	I0/I4056/net13	I0/I4056/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4062/T1	I0/I4062/net13	I0/I4062/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4064/T1	I0/I4064/net13	I0/I4064/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4053/T1	I0/I4053/net13	I0/I4053/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4067/T1	I0/I4067/net13	I0/I4067/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4061/T1	I0/I4061/net13	I0/I4061/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4065/T1	I0/I4065/net13	I0/I4065/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4046/T0	vdd	I0/I4046/net13	I0/I4046/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4047/T0	vdd	I0/I4047/net13	I0/I4047/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4054/T0	vdd	I0/I4054/net13	I0/I4054/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4056/T0	vdd	I0/I4056/net13	I0/I4056/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4062/T0	vdd	I0/I4062/net13	I0/I4062/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4064/T0	vdd	I0/I4064/net13	I0/I4064/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4053/T0	vdd	I0/I4053/net13	I0/I4053/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4067/T0	vdd	I0/I4067/net13	I0/I4067/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4061/T0	vdd	I0/I4061/net13	I0/I4061/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4065/T0	vdd	I0/I4065/net13	I0/I4065/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4142/T1	I0/I4142/net13	I0/I4142/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4143/T1	I0/I4143/net13	I0/I4143/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4150/T1	I0/I4150/net13	I0/I4150/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4152/T1	I0/I4152/net13	I0/I4152/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4158/T1	I0/I4158/net13	I0/I4158/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4160/T1	I0/I4160/net13	I0/I4160/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4149/T1	I0/I4149/net13	I0/I4149/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4163/T1	I0/I4163/net13	I0/I4163/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4157/T1	I0/I4157/net13	I0/I4157/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4161/T1	I0/I4161/net13	I0/I4161/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4142/T0	vdd	I0/I4142/net13	I0/I4142/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4143/T0	vdd	I0/I4143/net13	I0/I4143/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4150/T0	vdd	I0/I4150/net13	I0/I4150/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4152/T0	vdd	I0/I4152/net13	I0/I4152/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4158/T0	vdd	I0/I4158/net13	I0/I4158/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4160/T0	vdd	I0/I4160/net13	I0/I4160/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4149/T0	vdd	I0/I4149/net13	I0/I4149/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4163/T0	vdd	I0/I4163/net13	I0/I4163/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4157/T0	vdd	I0/I4157/net13	I0/I4157/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4161/T0	vdd	I0/I4161/net13	I0/I4161/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4174/T1	I0/I4174/net13	I0/I4174/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4175/T1	I0/I4175/net13	I0/I4175/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4182/T1	I0/I4182/net13	I0/I4182/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4184/T1	I0/I4184/net13	I0/I4184/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4190/T1	I0/I4190/net13	I0/I4190/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4192/T1	I0/I4192/net13	I0/I4192/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4181/T1	I0/I4181/net13	I0/I4181/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4195/T1	I0/I4195/net13	I0/I4195/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4189/T1	I0/I4189/net13	I0/I4189/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4193/T1	I0/I4193/net13	I0/I4193/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4174/T0	vdd	I0/I4174/net13	I0/I4174/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4175/T0	vdd	I0/I4175/net13	I0/I4175/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4182/T0	vdd	I0/I4182/net13	I0/I4182/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4184/T0	vdd	I0/I4184/net13	I0/I4184/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4190/T0	vdd	I0/I4190/net13	I0/I4190/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4192/T0	vdd	I0/I4192/net13	I0/I4192/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4181/T0	vdd	I0/I4181/net13	I0/I4181/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4195/T0	vdd	I0/I4195/net13	I0/I4195/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4189/T0	vdd	I0/I4189/net13	I0/I4189/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4193/T0	vdd	I0/I4193/net13	I0/I4193/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4206/T1	I0/I4206/net13	I0/I4206/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4207/T1	I0/I4207/net13	I0/I4207/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4214/T1	I0/I4214/net13	I0/I4214/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4216/T1	I0/I4216/net13	I0/I4216/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4222/T1	I0/I4222/net13	I0/I4222/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4224/T1	I0/I4224/net13	I0/I4224/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4213/T1	I0/I4213/net13	I0/I4213/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4227/T1	I0/I4227/net13	I0/I4227/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4221/T1	I0/I4221/net13	I0/I4221/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4225/T1	I0/I4225/net13	I0/I4225/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4077/T0	vdd	I0/I4077/net13	I0/I4077/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4063/T0	vdd	I0/I4063/net13	I0/I4063/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4074/T0	vdd	I0/I4074/net13	I0/I4074/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4073/T0	vdd	I0/I4073/net13	I0/I4073/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.4e-15 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4077/T1	I0/I4077/net13	I0/I4077/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4063/T1	I0/I4063/net13	I0/I4063/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4074/T1	I0/I4074/net13	I0/I4074/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4073/T1	I0/I4073/net13	I0/I4073/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.8e-15 panw8=3.08e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4173/T0	vdd	I0/I4173/net13	I0/I4173/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4159/T0	vdd	I0/I4159/net13	I0/I4159/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4170/T0	vdd	I0/I4170/net13	I0/I4170/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4169/T0	vdd	I0/I4169/net13	I0/I4169/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4173/T1	I0/I4173/net13	I0/I4173/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4159/T1	I0/I4159/net13	I0/I4159/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4170/T1	I0/I4170/net13	I0/I4170/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4169/T1	I0/I4169/net13	I0/I4169/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4205/T0	vdd	I0/I4205/net13	I0/I4205/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4191/T0	vdd	I0/I4191/net13	I0/I4191/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4202/T0	vdd	I0/I4202/net13	I0/I4202/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4201/T0	vdd	I0/I4201/net13	I0/I4201/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4205/T1	I0/I4205/net13	I0/I4205/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4191/T1	I0/I4191/net13	I0/I4191/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4202/T1	I0/I4202/net13	I0/I4202/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4201/T1	I0/I4201/net13	I0/I4201/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4237/T1	I0/I4237/net13	I0/I4237/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4223/T1	I0/I4223/net13	I0/I4223/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4234/T1	I0/I4234/net13	I0/I4234/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4233/T1	I0/I4233/net13	I0/I4233/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4210/T1	I0/I4210/net13	I0/I4210/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4178/T0	vdd	I0/I4178/net13	I0/I4178/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4178/T1	I0/I4178/net13	I0/I4178/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4146/T0	vdd	I0/I4146/net13	I0/I4146/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4146/T1	I0/I4146/net13	I0/I4146/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4050/T0	vdd	I0/I4050/net13	I0/I4050/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.36e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4050/T1	I0/I4050/net13	I0/I4050/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI109/T0	BL39	y4bar	p10	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI110/T0	p10bar	y3bar	BL38bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI111/T0	BL38	y3bar	p10	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI112/T0	p10bar	y2bar	BL37bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI113/T0	BL37	y2bar	p10	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI114/T0	p10bar	y1bar	BL36bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI115/T0	BL36	y1bar	p10	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=9.12e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T14	I32/net7	p9	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T15	p9bar	net681	I32/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T0	vdd	I11/net24	I11/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T1	I11/net20	I11/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T9	vdd	I11/net20	I11/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI11/T10	data9	I11/net8	vdd	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T10	I33/net23	data9	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T13	I33/net15	net681	p10	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T12	vdd	I33/net23	I33/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=3.06e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T14	I33/net7	p10	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.36e-13 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI33/T15	p10bar	net681	I33/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.64e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4206/T0	vdd	I0/I4206/net13	I0/I4206/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4207/T0	vdd	I0/I4207/net13	I0/I4207/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4214/T0	vdd	I0/I4214/net13	I0/I4214/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4216/T0	vdd	I0/I4216/net13	I0/I4216/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4222/T0	vdd	I0/I4222/net13	I0/I4222/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4224/T0	vdd	I0/I4224/net13	I0/I4224/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4213/T0	vdd	I0/I4213/net13	I0/I4213/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4227/T0	vdd	I0/I4227/net13	I0/I4227/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4221/T0	vdd	I0/I4221/net13	I0/I4221/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4225/T0	vdd	I0/I4225/net13	I0/I4225/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3918/T1	I0/I3918/net13	I0/I3918/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3919/T1	I0/I3919/net13	I0/I3919/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3926/T1	I0/I3926/net13	I0/I3926/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3928/T1	I0/I3928/net13	I0/I3928/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3934/T1	I0/I3934/net13	I0/I3934/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3936/T1	I0/I3936/net13	I0/I3936/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3925/T1	I0/I3925/net13	I0/I3925/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3939/T1	I0/I3939/net13	I0/I3939/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3933/T1	I0/I3933/net13	I0/I3933/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3937/T1	I0/I3937/net13	I0/I3937/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3918/T0	vdd	I0/I3918/net13	I0/I3918/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3919/T0	vdd	I0/I3919/net13	I0/I3919/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3926/T0	vdd	I0/I3926/net13	I0/I3926/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3928/T0	vdd	I0/I3928/net13	I0/I3928/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3934/T0	vdd	I0/I3934/net13	I0/I3934/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3936/T0	vdd	I0/I3936/net13	I0/I3936/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3925/T0	vdd	I0/I3925/net13	I0/I3925/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3939/T0	vdd	I0/I3939/net13	I0/I3939/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3933/T0	vdd	I0/I3933/net13	I0/I3933/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3937/T0	vdd	I0/I3937/net13	I0/I3937/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3950/T1	I0/I3950/net13	I0/I3950/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3951/T1	I0/I3951/net13	I0/I3951/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3958/T1	I0/I3958/net13	I0/I3958/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3960/T1	I0/I3960/net13	I0/I3960/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3966/T1	I0/I3966/net13	I0/I3966/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3968/T1	I0/I3968/net13	I0/I3968/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3957/T1	I0/I3957/net13	I0/I3957/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3971/T1	I0/I3971/net13	I0/I3971/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3965/T1	I0/I3965/net13	I0/I3965/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3969/T1	I0/I3969/net13	I0/I3969/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3950/T0	vdd	I0/I3950/net13	I0/I3950/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3951/T0	vdd	I0/I3951/net13	I0/I3951/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3958/T0	vdd	I0/I3958/net13	I0/I3958/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3960/T0	vdd	I0/I3960/net13	I0/I3960/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3966/T0	vdd	I0/I3966/net13	I0/I3966/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3968/T0	vdd	I0/I3968/net13	I0/I3968/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3957/T0	vdd	I0/I3957/net13	I0/I3957/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3971/T0	vdd	I0/I3971/net13	I0/I3971/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3965/T0	vdd	I0/I3965/net13	I0/I3965/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3969/T0	vdd	I0/I3969/net13	I0/I3969/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3982/T1	I0/I3982/net13	I0/I3982/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3983/T1	I0/I3983/net13	I0/I3983/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3990/T1	I0/I3990/net13	I0/I3990/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3992/T1	I0/I3992/net13	I0/I3992/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3998/T1	I0/I3998/net13	I0/I3998/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4000/T1	I0/I4000/net13	I0/I4000/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3989/T1	I0/I3989/net13	I0/I3989/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4003/T1	I0/I4003/net13	I0/I4003/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3997/T1	I0/I3997/net13	I0/I3997/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4001/T1	I0/I4001/net13	I0/I4001/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3982/T0	vdd	I0/I3982/net13	I0/I3982/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3983/T0	vdd	I0/I3983/net13	I0/I3983/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3990/T0	vdd	I0/I3990/net13	I0/I3990/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3992/T0	vdd	I0/I3992/net13	I0/I3992/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3998/T0	vdd	I0/I3998/net13	I0/I3998/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4000/T0	vdd	I0/I4000/net13	I0/I4000/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3989/T0	vdd	I0/I3989/net13	I0/I3989/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4003/T0	vdd	I0/I4003/net13	I0/I4003/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3997/T0	vdd	I0/I3997/net13	I0/I3997/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4001/T0	vdd	I0/I4001/net13	I0/I4001/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4237/T0	vdd	I0/I4237/net13	I0/I4237/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4223/T0	vdd	I0/I4223/net13	I0/I4223/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4234/T0	vdd	I0/I4234/net13	I0/I4234/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4233/T0	vdd	I0/I4233/net13	I0/I4233/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3949/T0	vdd	I0/I3949/net13	I0/I3949/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3935/T0	vdd	I0/I3935/net13	I0/I3935/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3946/T0	vdd	I0/I3946/net13	I0/I3946/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3945/T0	vdd	I0/I3945/net13	I0/I3945/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3949/T1	I0/I3949/net13	I0/I3949/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3935/T1	I0/I3935/net13	I0/I3935/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3946/T1	I0/I3946/net13	I0/I3946/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3945/T1	I0/I3945/net13	I0/I3945/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3981/T0	vdd	I0/I3981/net13	I0/I3981/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3967/T0	vdd	I0/I3967/net13	I0/I3967/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3978/T0	vdd	I0/I3978/net13	I0/I3978/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3977/T0	vdd	I0/I3977/net13	I0/I3977/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3981/T1	I0/I3981/net13	I0/I3981/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3967/T1	I0/I3967/net13	I0/I3967/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3978/T1	I0/I3978/net13	I0/I3978/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3977/T1	I0/I3977/net13	I0/I3977/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4013/T0	vdd	I0/I4013/net13	I0/I4013/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3999/T0	vdd	I0/I3999/net13	I0/I3999/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4010/T0	vdd	I0/I4010/net13	I0/I4010/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4009/T0	vdd	I0/I4009/net13	I0/I4009/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4013/T1	I0/I4013/net13	I0/I4013/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3999/T1	I0/I3999/net13	I0/I3999/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4010/T1	I0/I4010/net13	I0/I4010/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4009/T1	I0/I4009/net13	I0/I4009/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3986/T0	vdd	I0/I3986/net13	I0/I3986/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3986/T1	I0/I3986/net13	I0/I3986/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3954/T0	vdd	I0/I3954/net13	I0/I3954/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3954/T1	I0/I3954/net13	I0/I3954/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3922/T0	vdd	I0/I3922/net13	I0/I3922/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3922/T1	I0/I3922/net13	I0/I3922/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4210/T0	vdd	I0/I4210/net13	I0/I4210/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI102/T0	p9bar	y3bar	BL34bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI103/T0	BL34	y3bar	p9	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI104/T0	p9bar	y2bar	BL33bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI105/T0	BL33	y2bar	p9	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI106/T0	p9bar	y1bar	BL32bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI107/T0	BL32	y1bar	p9	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI108/T0	p10bar	y4bar	BL39bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T13	I31/net15	net681	p8	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T12	vdd	I31/net23	I31/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T14	I31/net7	p8	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T15	p8bar	net681	I31/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T0	vdd	I10/net24	I10/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T1	I10/net20	I10/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T9	vdd	I10/net20	I10/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI10/T10	data8	I10/net8	vdd	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T10	I32/net23	data8	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T13	I32/net15	net681	p9	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI32/T12	vdd	I32/net23	I32/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI147/T1	vdd	clkout	BL28bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3804/T0	vdd	I0/I3804/net13	I0/I3804/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI147/T2	BL28	clkout	BL28bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI147/T0	BL28	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3804/T1	I0/I3804/net13	I0/I3804/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI154/T1	vdd	clkout	BL35bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4028/T0	vdd	I0/I4028/net13	I0/I4028/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI154/T2	BL35	clkout	BL35bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI154/T0	BL35	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4028/T1	I0/I4028/net13	I0/I4028/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI149/T0	BL30	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3868/T1	I0/I3868/net13	I0/I3868/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI148/T1	vdd	clkout	BL29bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3836/T0	vdd	I0/I3836/net13	I0/I3836/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI148/T2	BL29	clkout	BL29bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI148/T0	BL29	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3836/T1	I0/I3836/net13	I0/I3836/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI149/T2	BL30	clkout	BL30bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI150/T1	vdd	clkout	BL31bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3900/T0	vdd	I0/I3900/net13	I0/I3900/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI150/T2	BL31	clkout	BL31bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI150/T0	BL31	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3900/T1	I0/I3900/net13	I0/I3900/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI149/T1	vdd	clkout	BL30bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3868/T0	vdd	I0/I3868/net13	I0/I3868/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI144/T1	vdd	clkout	BL25bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3708/T0	vdd	I0/I3708/net13	I0/I3708/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI144/T2	BL25	clkout	BL25bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI144/T0	BL25	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3708/T1	I0/I3708/net13	I0/I3708/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI143/T1	vdd	clkout	BL24bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3676/T0	vdd	I0/I3676/net13	I0/I3676/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI143/T2	BL24	clkout	BL24bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI143/T0	BL24	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3676/T1	I0/I3676/net13	I0/I3676/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3796/T0	vdd	I0/I3796/net13	I0/I3796/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3795/T0	vdd	I0/I3795/net13	I0/I3795/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3796/T1	I0/I3796/net13	I0/I3796/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3795/T1	I0/I3795/net13	I0/I3795/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4020/T0	vdd	I0/I4020/net13	I0/I4020/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4019/T0	vdd	I0/I4019/net13	I0/I4019/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4020/T1	I0/I4020/net13	I0/I4020/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4019/T1	I0/I4019/net13	I0/I4019/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3860/T1	I0/I3860/net13	I0/I3860/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3859/T1	I0/I3859/net13	I0/I3859/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3828/T0	vdd	I0/I3828/net13	I0/I3828/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3827/T0	vdd	I0/I3827/net13	I0/I3827/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3828/T1	I0/I3828/net13	I0/I3828/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3827/T1	I0/I3827/net13	I0/I3827/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3892/T0	vdd	I0/I3892/net13	I0/I3892/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3891/T0	vdd	I0/I3891/net13	I0/I3891/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3892/T1	I0/I3892/net13	I0/I3892/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3891/T1	I0/I3891/net13	I0/I3891/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3860/T0	vdd	I0/I3860/net13	I0/I3860/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3859/T0	vdd	I0/I3859/net13	I0/I3859/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3700/T0	vdd	I0/I3700/net13	I0/I3700/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3699/T0	vdd	I0/I3699/net13	I0/I3699/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3700/T1	I0/I3700/net13	I0/I3700/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3699/T1	I0/I3699/net13	I0/I3699/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3668/T0	vdd	I0/I3668/net13	I0/I3668/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3667/T0	vdd	I0/I3667/net13	I0/I3667/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3668/T1	I0/I3668/net13	I0/I3668/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3667/T1	I0/I3667/net13	I0/I3667/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4044/T0	vdd	I0/I4044/net13	I0/I4044/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4025/T0	vdd	I0/I4025/net13	I0/I4025/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4040/T0	vdd	I0/I4040/net13	I0/I4040/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4038/T0	vdd	I0/I4038/net13	I0/I4038/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4044/T1	I0/I4044/net13	I0/I4044/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4025/T1	I0/I4025/net13	I0/I4025/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4040/T1	I0/I4040/net13	I0/I4040/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4038/T1	I0/I4038/net13	I0/I4038/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3820/T0	vdd	I0/I3820/net13	I0/I3820/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3801/T0	vdd	I0/I3801/net13	I0/I3801/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3816/T0	vdd	I0/I3816/net13	I0/I3816/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3814/T0	vdd	I0/I3814/net13	I0/I3814/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3820/T1	I0/I3820/net13	I0/I3820/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3801/T1	I0/I3801/net13	I0/I3801/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3816/T1	I0/I3816/net13	I0/I3816/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3814/T1	I0/I3814/net13	I0/I3814/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3852/T0	vdd	I0/I3852/net13	I0/I3852/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3833/T0	vdd	I0/I3833/net13	I0/I3833/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3848/T0	vdd	I0/I3848/net13	I0/I3848/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3846/T0	vdd	I0/I3846/net13	I0/I3846/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3852/T1	I0/I3852/net13	I0/I3852/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3833/T1	I0/I3833/net13	I0/I3833/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3848/T1	I0/I3848/net13	I0/I3848/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3846/T1	I0/I3846/net13	I0/I3846/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3884/T1	I0/I3884/net13	I0/I3884/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3865/T1	I0/I3865/net13	I0/I3865/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3880/T1	I0/I3880/net13	I0/I3880/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3878/T1	I0/I3878/net13	I0/I3878/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3884/T0	vdd	I0/I3884/net13	I0/I3884/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3865/T0	vdd	I0/I3865/net13	I0/I3865/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3880/T0	vdd	I0/I3880/net13	I0/I3880/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3878/T0	vdd	I0/I3878/net13	I0/I3878/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3916/T0	vdd	I0/I3916/net13	I0/I3916/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3897/T0	vdd	I0/I3897/net13	I0/I3897/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3912/T0	vdd	I0/I3912/net13	I0/I3912/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3910/T0	vdd	I0/I3910/net13	I0/I3910/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3916/T1	I0/I3916/net13	I0/I3916/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3897/T1	I0/I3897/net13	I0/I3897/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3912/T1	I0/I3912/net13	I0/I3912/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3910/T1	I0/I3910/net13	I0/I3910/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3692/T0	vdd	I0/I3692/net13	I0/I3692/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3673/T0	vdd	I0/I3673/net13	I0/I3673/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3688/T0	vdd	I0/I3688/net13	I0/I3688/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3686/T0	vdd	I0/I3686/net13	I0/I3686/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3692/T1	I0/I3692/net13	I0/I3692/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3673/T1	I0/I3673/net13	I0/I3673/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3688/T1	I0/I3688/net13	I0/I3688/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3686/T1	I0/I3686/net13	I0/I3686/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3724/T0	vdd	I0/I3724/net13	I0/I3724/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3705/T0	vdd	I0/I3705/net13	I0/I3705/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3720/T0	vdd	I0/I3720/net13	I0/I3720/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3718/T0	vdd	I0/I3718/net13	I0/I3718/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3724/T1	I0/I3724/net13	I0/I3724/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3705/T1	I0/I3705/net13	I0/I3705/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3720/T1	I0/I3720/net13	I0/I3720/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3718/T1	I0/I3718/net13	I0/I3718/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4034/T1	I0/I4034/net13	I0/I4034/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4026/T1	I0/I4026/net13	I0/I4026/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4027/T1	I0/I4027/net13	I0/I4027/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4017/T1	I0/I4017/net13	I0/I4017/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4043/T1	I0/I4043/net13	I0/I4043/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4037/T1	I0/I4037/net13	I0/I4037/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4023/T1	I0/I4023/net13	I0/I4023/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4016/T1	I0/I4016/net13	I0/I4016/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4039/T1	I0/I4039/net13	I0/I4039/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4036/T1	I0/I4036/net13	I0/I4036/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4034/T0	vdd	I0/I4034/net13	I0/I4034/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4026/T0	vdd	I0/I4026/net13	I0/I4026/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4027/T0	vdd	I0/I4027/net13	I0/I4027/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4017/T0	vdd	I0/I4017/net13	I0/I4017/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4043/T0	vdd	I0/I4043/net13	I0/I4043/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4037/T0	vdd	I0/I4037/net13	I0/I4037/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4023/T0	vdd	I0/I4023/net13	I0/I4023/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4016/T0	vdd	I0/I4016/net13	I0/I4016/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4039/T0	vdd	I0/I4039/net13	I0/I4039/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4036/T0	vdd	I0/I4036/net13	I0/I4036/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3810/T1	I0/I3810/net13	I0/I3810/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3802/T1	I0/I3802/net13	I0/I3802/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3803/T1	I0/I3803/net13	I0/I3803/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3793/T1	I0/I3793/net13	I0/I3793/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3819/T1	I0/I3819/net13	I0/I3819/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3813/T1	I0/I3813/net13	I0/I3813/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3799/T1	I0/I3799/net13	I0/I3799/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3792/T1	I0/I3792/net13	I0/I3792/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3815/T1	I0/I3815/net13	I0/I3815/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3812/T1	I0/I3812/net13	I0/I3812/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3810/T0	vdd	I0/I3810/net13	I0/I3810/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3802/T0	vdd	I0/I3802/net13	I0/I3802/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3803/T0	vdd	I0/I3803/net13	I0/I3803/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3793/T0	vdd	I0/I3793/net13	I0/I3793/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3819/T0	vdd	I0/I3819/net13	I0/I3819/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3813/T0	vdd	I0/I3813/net13	I0/I3813/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3799/T0	vdd	I0/I3799/net13	I0/I3799/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3792/T0	vdd	I0/I3792/net13	I0/I3792/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3815/T0	vdd	I0/I3815/net13	I0/I3815/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3812/T0	vdd	I0/I3812/net13	I0/I3812/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3842/T1	I0/I3842/net13	I0/I3842/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3834/T1	I0/I3834/net13	I0/I3834/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3835/T1	I0/I3835/net13	I0/I3835/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3825/T1	I0/I3825/net13	I0/I3825/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3851/T1	I0/I3851/net13	I0/I3851/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3845/T1	I0/I3845/net13	I0/I3845/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3831/T1	I0/I3831/net13	I0/I3831/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3824/T1	I0/I3824/net13	I0/I3824/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3847/T1	I0/I3847/net13	I0/I3847/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3844/T1	I0/I3844/net13	I0/I3844/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3842/T0	vdd	I0/I3842/net13	I0/I3842/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3834/T0	vdd	I0/I3834/net13	I0/I3834/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3835/T0	vdd	I0/I3835/net13	I0/I3835/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3825/T0	vdd	I0/I3825/net13	I0/I3825/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3851/T0	vdd	I0/I3851/net13	I0/I3851/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3845/T0	vdd	I0/I3845/net13	I0/I3845/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3831/T0	vdd	I0/I3831/net13	I0/I3831/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3824/T0	vdd	I0/I3824/net13	I0/I3824/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3847/T0	vdd	I0/I3847/net13	I0/I3847/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3844/T0	vdd	I0/I3844/net13	I0/I3844/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3874/T1	I0/I3874/net13	I0/I3874/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3866/T1	I0/I3866/net13	I0/I3866/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3867/T1	I0/I3867/net13	I0/I3867/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3857/T1	I0/I3857/net13	I0/I3857/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3883/T1	I0/I3883/net13	I0/I3883/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3877/T1	I0/I3877/net13	I0/I3877/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3863/T1	I0/I3863/net13	I0/I3863/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3856/T1	I0/I3856/net13	I0/I3856/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3879/T1	I0/I3879/net13	I0/I3879/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3876/T1	I0/I3876/net13	I0/I3876/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3874/T0	vdd	I0/I3874/net13	I0/I3874/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3866/T0	vdd	I0/I3866/net13	I0/I3866/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3867/T0	vdd	I0/I3867/net13	I0/I3867/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3857/T0	vdd	I0/I3857/net13	I0/I3857/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3883/T0	vdd	I0/I3883/net13	I0/I3883/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3877/T0	vdd	I0/I3877/net13	I0/I3877/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3863/T0	vdd	I0/I3863/net13	I0/I3863/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3856/T0	vdd	I0/I3856/net13	I0/I3856/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3879/T0	vdd	I0/I3879/net13	I0/I3879/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3876/T0	vdd	I0/I3876/net13	I0/I3876/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3906/T1	I0/I3906/net13	I0/I3906/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3898/T1	I0/I3898/net13	I0/I3898/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3899/T1	I0/I3899/net13	I0/I3899/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3889/T1	I0/I3889/net13	I0/I3889/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3915/T1	I0/I3915/net13	I0/I3915/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3909/T1	I0/I3909/net13	I0/I3909/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3895/T1	I0/I3895/net13	I0/I3895/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3888/T1	I0/I3888/net13	I0/I3888/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3911/T1	I0/I3911/net13	I0/I3911/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3908/T1	I0/I3908/net13	I0/I3908/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3906/T0	vdd	I0/I3906/net13	I0/I3906/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3898/T0	vdd	I0/I3898/net13	I0/I3898/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3899/T0	vdd	I0/I3899/net13	I0/I3899/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3889/T0	vdd	I0/I3889/net13	I0/I3889/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3915/T0	vdd	I0/I3915/net13	I0/I3915/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3909/T0	vdd	I0/I3909/net13	I0/I3909/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3895/T0	vdd	I0/I3895/net13	I0/I3895/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3888/T0	vdd	I0/I3888/net13	I0/I3888/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3911/T0	vdd	I0/I3911/net13	I0/I3911/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3908/T0	vdd	I0/I3908/net13	I0/I3908/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3682/T1	I0/I3682/net13	I0/I3682/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3674/T1	I0/I3674/net13	I0/I3674/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3675/T1	I0/I3675/net13	I0/I3675/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3665/T1	I0/I3665/net13	I0/I3665/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3691/T1	I0/I3691/net13	I0/I3691/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3685/T1	I0/I3685/net13	I0/I3685/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3671/T1	I0/I3671/net13	I0/I3671/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3664/T1	I0/I3664/net13	I0/I3664/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3687/T1	I0/I3687/net13	I0/I3687/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3684/T1	I0/I3684/net13	I0/I3684/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3682/T0	vdd	I0/I3682/net13	I0/I3682/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3674/T0	vdd	I0/I3674/net13	I0/I3674/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3675/T0	vdd	I0/I3675/net13	I0/I3675/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3665/T0	vdd	I0/I3665/net13	I0/I3665/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3691/T0	vdd	I0/I3691/net13	I0/I3691/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3685/T0	vdd	I0/I3685/net13	I0/I3685/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3671/T0	vdd	I0/I3671/net13	I0/I3671/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3664/T0	vdd	I0/I3664/net13	I0/I3664/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3687/T0	vdd	I0/I3687/net13	I0/I3687/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3684/T0	vdd	I0/I3684/net13	I0/I3684/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3714/T1	I0/I3714/net13	I0/I3714/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3706/T1	I0/I3706/net13	I0/I3706/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3707/T1	I0/I3707/net13	I0/I3707/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3697/T1	I0/I3697/net13	I0/I3697/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3723/T1	I0/I3723/net13	I0/I3723/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3717/T1	I0/I3717/net13	I0/I3717/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3703/T1	I0/I3703/net13	I0/I3703/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3696/T1	I0/I3696/net13	I0/I3696/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3719/T1	I0/I3719/net13	I0/I3719/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3716/T1	I0/I3716/net13	I0/I3716/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3714/T0	vdd	I0/I3714/net13	I0/I3714/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3706/T0	vdd	I0/I3706/net13	I0/I3706/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3707/T0	vdd	I0/I3707/net13	I0/I3707/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3697/T0	vdd	I0/I3697/net13	I0/I3697/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3723/T0	vdd	I0/I3723/net13	I0/I3723/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3717/T0	vdd	I0/I3717/net13	I0/I3717/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3703/T0	vdd	I0/I3703/net13	I0/I3703/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3696/T0	vdd	I0/I3696/net13	I0/I3696/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3719/T0	vdd	I0/I3719/net13	I0/I3719/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3716/T0	vdd	I0/I3716/net13	I0/I3716/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4014/T1	I0/I4014/net13	I0/I4014/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4015/T1	I0/I4015/net13	I0/I4015/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4022/T1	I0/I4022/net13	I0/I4022/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4024/T1	I0/I4024/net13	I0/I4024/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4030/T1	I0/I4030/net13	I0/I4030/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4032/T1	I0/I4032/net13	I0/I4032/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4021/T1	I0/I4021/net13	I0/I4021/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4035/T1	I0/I4035/net13	I0/I4035/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4029/T1	I0/I4029/net13	I0/I4029/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4033/T1	I0/I4033/net13	I0/I4033/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4014/T0	vdd	I0/I4014/net13	I0/I4014/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4015/T0	vdd	I0/I4015/net13	I0/I4015/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4022/T0	vdd	I0/I4022/net13	I0/I4022/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4024/T0	vdd	I0/I4024/net13	I0/I4024/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4030/T0	vdd	I0/I4030/net13	I0/I4030/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4032/T0	vdd	I0/I4032/net13	I0/I4032/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4021/T0	vdd	I0/I4021/net13	I0/I4021/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4035/T0	vdd	I0/I4035/net13	I0/I4035/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4029/T0	vdd	I0/I4029/net13	I0/I4029/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4033/T0	vdd	I0/I4033/net13	I0/I4033/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3790/T1	I0/I3790/net13	I0/I3790/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3791/T1	I0/I3791/net13	I0/I3791/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3798/T1	I0/I3798/net13	I0/I3798/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3800/T1	I0/I3800/net13	I0/I3800/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3806/T1	I0/I3806/net13	I0/I3806/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3808/T1	I0/I3808/net13	I0/I3808/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3797/T1	I0/I3797/net13	I0/I3797/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3811/T1	I0/I3811/net13	I0/I3811/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3805/T1	I0/I3805/net13	I0/I3805/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3809/T1	I0/I3809/net13	I0/I3809/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3790/T0	vdd	I0/I3790/net13	I0/I3790/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3791/T0	vdd	I0/I3791/net13	I0/I3791/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3798/T0	vdd	I0/I3798/net13	I0/I3798/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3800/T0	vdd	I0/I3800/net13	I0/I3800/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3806/T0	vdd	I0/I3806/net13	I0/I3806/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3808/T0	vdd	I0/I3808/net13	I0/I3808/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3797/T0	vdd	I0/I3797/net13	I0/I3797/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3811/T0	vdd	I0/I3811/net13	I0/I3811/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3805/T0	vdd	I0/I3805/net13	I0/I3805/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3809/T0	vdd	I0/I3809/net13	I0/I3809/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3822/T1	I0/I3822/net13	I0/I3822/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3823/T1	I0/I3823/net13	I0/I3823/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3830/T1	I0/I3830/net13	I0/I3830/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3832/T1	I0/I3832/net13	I0/I3832/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3838/T1	I0/I3838/net13	I0/I3838/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3840/T1	I0/I3840/net13	I0/I3840/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3829/T1	I0/I3829/net13	I0/I3829/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3843/T1	I0/I3843/net13	I0/I3843/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3837/T1	I0/I3837/net13	I0/I3837/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3841/T1	I0/I3841/net13	I0/I3841/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3822/T0	vdd	I0/I3822/net13	I0/I3822/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3823/T0	vdd	I0/I3823/net13	I0/I3823/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3830/T0	vdd	I0/I3830/net13	I0/I3830/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3832/T0	vdd	I0/I3832/net13	I0/I3832/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3838/T0	vdd	I0/I3838/net13	I0/I3838/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3840/T0	vdd	I0/I3840/net13	I0/I3840/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3829/T0	vdd	I0/I3829/net13	I0/I3829/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3843/T0	vdd	I0/I3843/net13	I0/I3843/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3837/T0	vdd	I0/I3837/net13	I0/I3837/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3841/T0	vdd	I0/I3841/net13	I0/I3841/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3854/T1	I0/I3854/net13	I0/I3854/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3855/T1	I0/I3855/net13	I0/I3855/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3862/T1	I0/I3862/net13	I0/I3862/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3864/T1	I0/I3864/net13	I0/I3864/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3870/T1	I0/I3870/net13	I0/I3870/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3872/T1	I0/I3872/net13	I0/I3872/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3861/T1	I0/I3861/net13	I0/I3861/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3875/T1	I0/I3875/net13	I0/I3875/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3869/T1	I0/I3869/net13	I0/I3869/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3873/T1	I0/I3873/net13	I0/I3873/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4045/T0	vdd	I0/I4045/net13	I0/I4045/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4031/T0	vdd	I0/I4031/net13	I0/I4031/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4042/T0	vdd	I0/I4042/net13	I0/I4042/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4041/T0	vdd	I0/I4041/net13	I0/I4041/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4045/T1	I0/I4045/net13	I0/I4045/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4031/T1	I0/I4031/net13	I0/I4031/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4042/T1	I0/I4042/net13	I0/I4042/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4041/T1	I0/I4041/net13	I0/I4041/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3821/T0	vdd	I0/I3821/net13	I0/I3821/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3807/T0	vdd	I0/I3807/net13	I0/I3807/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3818/T0	vdd	I0/I3818/net13	I0/I3818/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3817/T0	vdd	I0/I3817/net13	I0/I3817/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3821/T1	I0/I3821/net13	I0/I3821/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3807/T1	I0/I3807/net13	I0/I3807/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3818/T1	I0/I3818/net13	I0/I3818/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3817/T1	I0/I3817/net13	I0/I3817/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3853/T0	vdd	I0/I3853/net13	I0/I3853/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3839/T0	vdd	I0/I3839/net13	I0/I3839/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3850/T0	vdd	I0/I3850/net13	I0/I3850/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3849/T0	vdd	I0/I3849/net13	I0/I3849/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3853/T1	I0/I3853/net13	I0/I3853/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3839/T1	I0/I3839/net13	I0/I3839/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3850/T1	I0/I3850/net13	I0/I3850/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3849/T1	I0/I3849/net13	I0/I3849/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3885/T1	I0/I3885/net13	I0/I3885/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3871/T1	I0/I3871/net13	I0/I3871/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3882/T1	I0/I3882/net13	I0/I3882/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3881/T1	I0/I3881/net13	I0/I3881/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3858/T1	I0/I3858/net13	I0/I3858/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3826/T0	vdd	I0/I3826/net13	I0/I3826/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3826/T1	I0/I3826/net13	I0/I3826/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3794/T0	vdd	I0/I3794/net13	I0/I3794/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3794/T1	I0/I3794/net13	I0/I3794/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4018/T0	vdd	I0/I4018/net13	I0/I4018/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I4018/T1	I0/I4018/net13	I0/I4018/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI95/T0	BL30	y3bar	p8	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI96/T0	p8bar	y2bar	BL29bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI97/T0	BL29	y2bar	p8	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI98/T0	p8bar	y1bar	BL28bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI99/T0	BL28	y1bar	p8	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI100/T0	p9bar	y4bar	BL35bar	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI101/T0	BL35	y4bar	p9	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T10	I29/net23	data6	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T13	I29/net15	net681	p7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T12	vdd	I29/net23	I29/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T14	I29/net7	p7	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI29/T15	p7bar	net681	I29/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T0	vdd	I8/net24	I8/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T1	I8/net20	I8/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T9	vdd	I8/net20	I8/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI8/T10	data7	I8/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI31/T10	I31/net23	data7	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3854/T0	vdd	I0/I3854/net13	I0/I3854/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3855/T0	vdd	I0/I3855/net13	I0/I3855/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3862/T0	vdd	I0/I3862/net13	I0/I3862/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3864/T0	vdd	I0/I3864/net13	I0/I3864/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3870/T0	vdd	I0/I3870/net13	I0/I3870/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3872/T0	vdd	I0/I3872/net13	I0/I3872/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3861/T0	vdd	I0/I3861/net13	I0/I3861/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3875/T0	vdd	I0/I3875/net13	I0/I3875/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3869/T0	vdd	I0/I3869/net13	I0/I3869/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3873/T0	vdd	I0/I3873/net13	I0/I3873/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3886/T1	I0/I3886/net13	I0/I3886/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3887/T1	I0/I3887/net13	I0/I3887/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3894/T1	I0/I3894/net13	I0/I3894/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3896/T1	I0/I3896/net13	I0/I3896/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3902/T1	I0/I3902/net13	I0/I3902/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3904/T1	I0/I3904/net13	I0/I3904/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3893/T1	I0/I3893/net13	I0/I3893/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3907/T1	I0/I3907/net13	I0/I3907/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3901/T1	I0/I3901/net13	I0/I3901/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3905/T1	I0/I3905/net13	I0/I3905/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3886/T0	vdd	I0/I3886/net13	I0/I3886/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3887/T0	vdd	I0/I3887/net13	I0/I3887/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3894/T0	vdd	I0/I3894/net13	I0/I3894/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3896/T0	vdd	I0/I3896/net13	I0/I3896/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3902/T0	vdd	I0/I3902/net13	I0/I3902/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3904/T0	vdd	I0/I3904/net13	I0/I3904/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3893/T0	vdd	I0/I3893/net13	I0/I3893/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3907/T0	vdd	I0/I3907/net13	I0/I3907/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3901/T0	vdd	I0/I3901/net13	I0/I3901/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3905/T0	vdd	I0/I3905/net13	I0/I3905/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3662/T1	I0/I3662/net13	I0/I3662/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3663/T1	I0/I3663/net13	I0/I3663/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3670/T1	I0/I3670/net13	I0/I3670/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3672/T1	I0/I3672/net13	I0/I3672/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3678/T1	I0/I3678/net13	I0/I3678/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3680/T1	I0/I3680/net13	I0/I3680/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3669/T1	I0/I3669/net13	I0/I3669/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3683/T1	I0/I3683/net13	I0/I3683/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3677/T1	I0/I3677/net13	I0/I3677/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3681/T1	I0/I3681/net13	I0/I3681/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3662/T0	vdd	I0/I3662/net13	I0/I3662/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3663/T0	vdd	I0/I3663/net13	I0/I3663/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3670/T0	vdd	I0/I3670/net13	I0/I3670/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3672/T0	vdd	I0/I3672/net13	I0/I3672/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3678/T0	vdd	I0/I3678/net13	I0/I3678/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3680/T0	vdd	I0/I3680/net13	I0/I3680/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3669/T0	vdd	I0/I3669/net13	I0/I3669/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3683/T0	vdd	I0/I3683/net13	I0/I3683/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3677/T0	vdd	I0/I3677/net13	I0/I3677/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3681/T0	vdd	I0/I3681/net13	I0/I3681/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3694/T1	I0/I3694/net13	I0/I3694/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3695/T1	I0/I3695/net13	I0/I3695/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3702/T1	I0/I3702/net13	I0/I3702/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3704/T1	I0/I3704/net13	I0/I3704/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3710/T1	I0/I3710/net13	I0/I3710/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3712/T1	I0/I3712/net13	I0/I3712/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3701/T1	I0/I3701/net13	I0/I3701/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3715/T1	I0/I3715/net13	I0/I3715/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3709/T1	I0/I3709/net13	I0/I3709/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3713/T1	I0/I3713/net13	I0/I3713/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3694/T0	vdd	I0/I3694/net13	I0/I3694/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3695/T0	vdd	I0/I3695/net13	I0/I3695/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3702/T0	vdd	I0/I3702/net13	I0/I3702/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3704/T0	vdd	I0/I3704/net13	I0/I3704/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3710/T0	vdd	I0/I3710/net13	I0/I3710/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3712/T0	vdd	I0/I3712/net13	I0/I3712/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3701/T0	vdd	I0/I3701/net13	I0/I3701/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3715/T0	vdd	I0/I3715/net13	I0/I3715/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3709/T0	vdd	I0/I3709/net13	I0/I3709/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3713/T0	vdd	I0/I3713/net13	I0/I3713/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3885/T0	vdd	I0/I3885/net13	I0/I3885/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3871/T0	vdd	I0/I3871/net13	I0/I3871/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3882/T0	vdd	I0/I3882/net13	I0/I3882/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3881/T0	vdd	I0/I3881/net13	I0/I3881/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3917/T0	vdd	I0/I3917/net13	I0/I3917/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3903/T0	vdd	I0/I3903/net13	I0/I3903/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3914/T0	vdd	I0/I3914/net13	I0/I3914/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3913/T0	vdd	I0/I3913/net13	I0/I3913/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3917/T1	I0/I3917/net13	I0/I3917/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3903/T1	I0/I3903/net13	I0/I3903/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3914/T1	I0/I3914/net13	I0/I3914/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3913/T1	I0/I3913/net13	I0/I3913/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3693/T0	vdd	I0/I3693/net13	I0/I3693/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3679/T0	vdd	I0/I3679/net13	I0/I3679/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3690/T0	vdd	I0/I3690/net13	I0/I3690/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3689/T0	vdd	I0/I3689/net13	I0/I3689/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3693/T1	I0/I3693/net13	I0/I3693/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3679/T1	I0/I3679/net13	I0/I3679/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3690/T1	I0/I3690/net13	I0/I3690/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3689/T1	I0/I3689/net13	I0/I3689/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3725/T0	vdd	I0/I3725/net13	I0/I3725/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3711/T0	vdd	I0/I3711/net13	I0/I3711/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3722/T0	vdd	I0/I3722/net13	I0/I3722/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3721/T0	vdd	I0/I3721/net13	I0/I3721/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3725/T1	I0/I3725/net13	I0/I3725/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3711/T1	I0/I3711/net13	I0/I3711/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3722/T1	I0/I3722/net13	I0/I3722/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3721/T1	I0/I3721/net13	I0/I3721/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3698/T0	vdd	I0/I3698/net13	I0/I3698/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3698/T1	I0/I3698/net13	I0/I3698/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3666/T0	vdd	I0/I3666/net13	I0/I3666/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3666/T1	I0/I3666/net13	I0/I3666/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3890/T0	vdd	I0/I3890/net13	I0/I3890/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3890/T1	I0/I3890/net13	I0/I3890/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3858/T0	vdd	I0/I3858/net13	I0/I3858/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI88/T0	p7bar	y2bar	BL25bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI89/T0	BL25	y2bar	p7	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI90/T0	p7bar	y1bar	BL24bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI91/T0	BL24	y1bar	p7	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI92/T0	p8bar	y4bar	BL31bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI93/T0	BL31	y4bar	p8	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI94/T0	p8bar	y3bar	BL30bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T9	vdd	I6/net20	I6/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T10	data5	I6/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T10	I28/net23	data5	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T13	I28/net15	net681	p6	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T12	vdd	I28/net23	I28/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T14	I28/net7	p6	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI28/T15	p6bar	net681	I28/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T0	vdd	I7/net24	I7/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T1	I7/net20	I7/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T9	vdd	I7/net20	I7/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI7/T10	data6	I7/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI87/T0	BL26	y3bar	p7	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI146/T1	vdd	clkout	BL27bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3772/T0	vdd	I0/I3772/net13	I0/I3772/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI146/T2	BL27	clkout	BL27bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI146/T0	BL27	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3772/T1	I0/I3772/net13	I0/I3772/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI145/T1	vdd	clkout	BL26bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3740/T0	vdd	I0/I3740/net13	I0/I3740/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI145/T2	BL26	clkout	BL26bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI145/T0	BL26	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3740/T1	I0/I3740/net13	I0/I3740/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI140/T0	BL21	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3580/T1	I0/I3580/net13	I0/I3580/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI139/T1	vdd	clkout	BL20bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3548/T0	vdd	I0/I3548/net13	I0/I3548/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI139/T2	BL20	clkout	BL20bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI139/T0	BL20	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3548/T1	I0/I3548/net13	I0/I3548/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI140/T2	BL21	clkout	BL21bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI141/T1	vdd	clkout	BL22bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3612/T0	vdd	I0/I3612/net13	I0/I3612/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI141/T2	BL22	clkout	BL22bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI141/T0	BL22	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3612/T1	I0/I3612/net13	I0/I3612/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI140/T1	vdd	clkout	BL21bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3580/T0	vdd	I0/I3580/net13	I0/I3580/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI135/T1	vdd	clkout	BL16bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3420/T0	vdd	I0/I3420/net13	I0/I3420/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI135/T2	BL16	clkout	BL16bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI135/T0	BL16	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3420/T1	I0/I3420/net13	I0/I3420/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI142/T1	vdd	clkout	BL23bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3644/T0	vdd	I0/I3644/net13	I0/I3644/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI142/T2	BL23	clkout	BL23bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI142/T0	BL23	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3644/T1	I0/I3644/net13	I0/I3644/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3764/T0	vdd	I0/I3764/net13	I0/I3764/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3763/T0	vdd	I0/I3763/net13	I0/I3763/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3764/T1	I0/I3764/net13	I0/I3764/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3763/T1	I0/I3763/net13	I0/I3763/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3732/T0	vdd	I0/I3732/net13	I0/I3732/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3731/T0	vdd	I0/I3731/net13	I0/I3731/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3732/T1	I0/I3732/net13	I0/I3732/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3731/T1	I0/I3731/net13	I0/I3731/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3572/T1	I0/I3572/net13	I0/I3572/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3571/T1	I0/I3571/net13	I0/I3571/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3540/T0	vdd	I0/I3540/net13	I0/I3540/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3539/T0	vdd	I0/I3539/net13	I0/I3539/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3540/T1	I0/I3540/net13	I0/I3540/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3539/T1	I0/I3539/net13	I0/I3539/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3604/T0	vdd	I0/I3604/net13	I0/I3604/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3603/T0	vdd	I0/I3603/net13	I0/I3603/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3604/T1	I0/I3604/net13	I0/I3604/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3603/T1	I0/I3603/net13	I0/I3603/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3572/T0	vdd	I0/I3572/net13	I0/I3572/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3571/T0	vdd	I0/I3571/net13	I0/I3571/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3412/T0	vdd	I0/I3412/net13	I0/I3412/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3411/T0	vdd	I0/I3411/net13	I0/I3411/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3412/T1	I0/I3412/net13	I0/I3412/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3411/T1	I0/I3411/net13	I0/I3411/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3636/T0	vdd	I0/I3636/net13	I0/I3636/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3635/T0	vdd	I0/I3635/net13	I0/I3635/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3636/T1	I0/I3636/net13	I0/I3636/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3635/T1	I0/I3635/net13	I0/I3635/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3756/T0	vdd	I0/I3756/net13	I0/I3756/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3737/T0	vdd	I0/I3737/net13	I0/I3737/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3752/T0	vdd	I0/I3752/net13	I0/I3752/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3750/T0	vdd	I0/I3750/net13	I0/I3750/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3756/T1	I0/I3756/net13	I0/I3756/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3737/T1	I0/I3737/net13	I0/I3737/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3752/T1	I0/I3752/net13	I0/I3752/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3750/T1	I0/I3750/net13	I0/I3750/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3788/T0	vdd	I0/I3788/net13	I0/I3788/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3769/T0	vdd	I0/I3769/net13	I0/I3769/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3784/T0	vdd	I0/I3784/net13	I0/I3784/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3782/T0	vdd	I0/I3782/net13	I0/I3782/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3788/T1	I0/I3788/net13	I0/I3788/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3769/T1	I0/I3769/net13	I0/I3769/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3784/T1	I0/I3784/net13	I0/I3784/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3782/T1	I0/I3782/net13	I0/I3782/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3564/T0	vdd	I0/I3564/net13	I0/I3564/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3545/T0	vdd	I0/I3545/net13	I0/I3545/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3560/T0	vdd	I0/I3560/net13	I0/I3560/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3558/T0	vdd	I0/I3558/net13	I0/I3558/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3564/T1	I0/I3564/net13	I0/I3564/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3545/T1	I0/I3545/net13	I0/I3545/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3560/T1	I0/I3560/net13	I0/I3560/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3558/T1	I0/I3558/net13	I0/I3558/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3596/T1	I0/I3596/net13	I0/I3596/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3577/T1	I0/I3577/net13	I0/I3577/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3592/T1	I0/I3592/net13	I0/I3592/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3590/T1	I0/I3590/net13	I0/I3590/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3596/T0	vdd	I0/I3596/net13	I0/I3596/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3577/T0	vdd	I0/I3577/net13	I0/I3577/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3592/T0	vdd	I0/I3592/net13	I0/I3592/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3590/T0	vdd	I0/I3590/net13	I0/I3590/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3628/T0	vdd	I0/I3628/net13	I0/I3628/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3609/T0	vdd	I0/I3609/net13	I0/I3609/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3624/T0	vdd	I0/I3624/net13	I0/I3624/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3622/T0	vdd	I0/I3622/net13	I0/I3622/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3628/T1	I0/I3628/net13	I0/I3628/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3609/T1	I0/I3609/net13	I0/I3609/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3624/T1	I0/I3624/net13	I0/I3624/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3622/T1	I0/I3622/net13	I0/I3622/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3660/T0	vdd	I0/I3660/net13	I0/I3660/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3641/T0	vdd	I0/I3641/net13	I0/I3641/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3656/T0	vdd	I0/I3656/net13	I0/I3656/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3654/T0	vdd	I0/I3654/net13	I0/I3654/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3660/T1	I0/I3660/net13	I0/I3660/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3641/T1	I0/I3641/net13	I0/I3641/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3656/T1	I0/I3656/net13	I0/I3656/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3654/T1	I0/I3654/net13	I0/I3654/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3436/T0	vdd	I0/I3436/net13	I0/I3436/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3417/T0	vdd	I0/I3417/net13	I0/I3417/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3432/T0	vdd	I0/I3432/net13	I0/I3432/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3430/T0	vdd	I0/I3430/net13	I0/I3430/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3436/T1	I0/I3436/net13	I0/I3436/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3417/T1	I0/I3417/net13	I0/I3417/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3432/T1	I0/I3432/net13	I0/I3432/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3430/T1	I0/I3430/net13	I0/I3430/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3746/T1	I0/I3746/net13	I0/I3746/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3738/T1	I0/I3738/net13	I0/I3738/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3739/T1	I0/I3739/net13	I0/I3739/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3729/T1	I0/I3729/net13	I0/I3729/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3755/T1	I0/I3755/net13	I0/I3755/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3749/T1	I0/I3749/net13	I0/I3749/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3735/T1	I0/I3735/net13	I0/I3735/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3728/T1	I0/I3728/net13	I0/I3728/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3751/T1	I0/I3751/net13	I0/I3751/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3748/T1	I0/I3748/net13	I0/I3748/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3746/T0	vdd	I0/I3746/net13	I0/I3746/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3738/T0	vdd	I0/I3738/net13	I0/I3738/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3739/T0	vdd	I0/I3739/net13	I0/I3739/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3729/T0	vdd	I0/I3729/net13	I0/I3729/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3755/T0	vdd	I0/I3755/net13	I0/I3755/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3749/T0	vdd	I0/I3749/net13	I0/I3749/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3735/T0	vdd	I0/I3735/net13	I0/I3735/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3728/T0	vdd	I0/I3728/net13	I0/I3728/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3751/T0	vdd	I0/I3751/net13	I0/I3751/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3748/T0	vdd	I0/I3748/net13	I0/I3748/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3778/T1	I0/I3778/net13	I0/I3778/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3770/T1	I0/I3770/net13	I0/I3770/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3771/T1	I0/I3771/net13	I0/I3771/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3761/T1	I0/I3761/net13	I0/I3761/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3787/T1	I0/I3787/net13	I0/I3787/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3781/T1	I0/I3781/net13	I0/I3781/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3767/T1	I0/I3767/net13	I0/I3767/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3760/T1	I0/I3760/net13	I0/I3760/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3783/T1	I0/I3783/net13	I0/I3783/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3780/T1	I0/I3780/net13	I0/I3780/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3778/T0	vdd	I0/I3778/net13	I0/I3778/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3770/T0	vdd	I0/I3770/net13	I0/I3770/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3771/T0	vdd	I0/I3771/net13	I0/I3771/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3761/T0	vdd	I0/I3761/net13	I0/I3761/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3787/T0	vdd	I0/I3787/net13	I0/I3787/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3781/T0	vdd	I0/I3781/net13	I0/I3781/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3767/T0	vdd	I0/I3767/net13	I0/I3767/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3760/T0	vdd	I0/I3760/net13	I0/I3760/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3783/T0	vdd	I0/I3783/net13	I0/I3783/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3780/T0	vdd	I0/I3780/net13	I0/I3780/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3554/T1	I0/I3554/net13	I0/I3554/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3546/T1	I0/I3546/net13	I0/I3546/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3547/T1	I0/I3547/net13	I0/I3547/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3537/T1	I0/I3537/net13	I0/I3537/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3563/T1	I0/I3563/net13	I0/I3563/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3557/T1	I0/I3557/net13	I0/I3557/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3543/T1	I0/I3543/net13	I0/I3543/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3536/T1	I0/I3536/net13	I0/I3536/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3559/T1	I0/I3559/net13	I0/I3559/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3556/T1	I0/I3556/net13	I0/I3556/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3554/T0	vdd	I0/I3554/net13	I0/I3554/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3546/T0	vdd	I0/I3546/net13	I0/I3546/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3547/T0	vdd	I0/I3547/net13	I0/I3547/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3537/T0	vdd	I0/I3537/net13	I0/I3537/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3563/T0	vdd	I0/I3563/net13	I0/I3563/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3557/T0	vdd	I0/I3557/net13	I0/I3557/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3543/T0	vdd	I0/I3543/net13	I0/I3543/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3536/T0	vdd	I0/I3536/net13	I0/I3536/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3559/T0	vdd	I0/I3559/net13	I0/I3559/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3556/T0	vdd	I0/I3556/net13	I0/I3556/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3586/T1	I0/I3586/net13	I0/I3586/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3578/T1	I0/I3578/net13	I0/I3578/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3579/T1	I0/I3579/net13	I0/I3579/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3569/T1	I0/I3569/net13	I0/I3569/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3595/T1	I0/I3595/net13	I0/I3595/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3589/T1	I0/I3589/net13	I0/I3589/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3575/T1	I0/I3575/net13	I0/I3575/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3568/T1	I0/I3568/net13	I0/I3568/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3591/T1	I0/I3591/net13	I0/I3591/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3588/T1	I0/I3588/net13	I0/I3588/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3586/T0	vdd	I0/I3586/net13	I0/I3586/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3578/T0	vdd	I0/I3578/net13	I0/I3578/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3579/T0	vdd	I0/I3579/net13	I0/I3579/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3569/T0	vdd	I0/I3569/net13	I0/I3569/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3595/T0	vdd	I0/I3595/net13	I0/I3595/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3589/T0	vdd	I0/I3589/net13	I0/I3589/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3575/T0	vdd	I0/I3575/net13	I0/I3575/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3568/T0	vdd	I0/I3568/net13	I0/I3568/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3591/T0	vdd	I0/I3591/net13	I0/I3591/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3588/T0	vdd	I0/I3588/net13	I0/I3588/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3618/T1	I0/I3618/net13	I0/I3618/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3610/T1	I0/I3610/net13	I0/I3610/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3611/T1	I0/I3611/net13	I0/I3611/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3601/T1	I0/I3601/net13	I0/I3601/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3627/T1	I0/I3627/net13	I0/I3627/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3621/T1	I0/I3621/net13	I0/I3621/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3607/T1	I0/I3607/net13	I0/I3607/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3600/T1	I0/I3600/net13	I0/I3600/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3623/T1	I0/I3623/net13	I0/I3623/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3620/T1	I0/I3620/net13	I0/I3620/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3618/T0	vdd	I0/I3618/net13	I0/I3618/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3610/T0	vdd	I0/I3610/net13	I0/I3610/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3611/T0	vdd	I0/I3611/net13	I0/I3611/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3601/T0	vdd	I0/I3601/net13	I0/I3601/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3627/T0	vdd	I0/I3627/net13	I0/I3627/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3621/T0	vdd	I0/I3621/net13	I0/I3621/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3607/T0	vdd	I0/I3607/net13	I0/I3607/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3600/T0	vdd	I0/I3600/net13	I0/I3600/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3623/T0	vdd	I0/I3623/net13	I0/I3623/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3620/T0	vdd	I0/I3620/net13	I0/I3620/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3650/T1	I0/I3650/net13	I0/I3650/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3642/T1	I0/I3642/net13	I0/I3642/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3643/T1	I0/I3643/net13	I0/I3643/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3633/T1	I0/I3633/net13	I0/I3633/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3659/T1	I0/I3659/net13	I0/I3659/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3653/T1	I0/I3653/net13	I0/I3653/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3639/T1	I0/I3639/net13	I0/I3639/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3632/T1	I0/I3632/net13	I0/I3632/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3655/T1	I0/I3655/net13	I0/I3655/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3652/T1	I0/I3652/net13	I0/I3652/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3650/T0	vdd	I0/I3650/net13	I0/I3650/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3642/T0	vdd	I0/I3642/net13	I0/I3642/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3643/T0	vdd	I0/I3643/net13	I0/I3643/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3633/T0	vdd	I0/I3633/net13	I0/I3633/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3659/T0	vdd	I0/I3659/net13	I0/I3659/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3653/T0	vdd	I0/I3653/net13	I0/I3653/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3639/T0	vdd	I0/I3639/net13	I0/I3639/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3632/T0	vdd	I0/I3632/net13	I0/I3632/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3655/T0	vdd	I0/I3655/net13	I0/I3655/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3652/T0	vdd	I0/I3652/net13	I0/I3652/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3426/T1	I0/I3426/net13	I0/I3426/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3418/T1	I0/I3418/net13	I0/I3418/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3419/T1	I0/I3419/net13	I0/I3419/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3409/T1	I0/I3409/net13	I0/I3409/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3435/T1	I0/I3435/net13	I0/I3435/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3429/T1	I0/I3429/net13	I0/I3429/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3415/T1	I0/I3415/net13	I0/I3415/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3408/T1	I0/I3408/net13	I0/I3408/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3431/T1	I0/I3431/net13	I0/I3431/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3428/T1	I0/I3428/net13	I0/I3428/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3426/T0	vdd	I0/I3426/net13	I0/I3426/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3418/T0	vdd	I0/I3418/net13	I0/I3418/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3419/T0	vdd	I0/I3419/net13	I0/I3419/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3409/T0	vdd	I0/I3409/net13	I0/I3409/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3435/T0	vdd	I0/I3435/net13	I0/I3435/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3429/T0	vdd	I0/I3429/net13	I0/I3429/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3415/T0	vdd	I0/I3415/net13	I0/I3415/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3408/T0	vdd	I0/I3408/net13	I0/I3408/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3431/T0	vdd	I0/I3431/net13	I0/I3431/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3428/T0	vdd	I0/I3428/net13	I0/I3428/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3726/T1	I0/I3726/net13	I0/I3726/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3727/T1	I0/I3727/net13	I0/I3727/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3734/T1	I0/I3734/net13	I0/I3734/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3736/T1	I0/I3736/net13	I0/I3736/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3742/T1	I0/I3742/net13	I0/I3742/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3744/T1	I0/I3744/net13	I0/I3744/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3733/T1	I0/I3733/net13	I0/I3733/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3747/T1	I0/I3747/net13	I0/I3747/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3741/T1	I0/I3741/net13	I0/I3741/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3745/T1	I0/I3745/net13	I0/I3745/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3726/T0	vdd	I0/I3726/net13	I0/I3726/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3727/T0	vdd	I0/I3727/net13	I0/I3727/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3734/T0	vdd	I0/I3734/net13	I0/I3734/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3736/T0	vdd	I0/I3736/net13	I0/I3736/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3742/T0	vdd	I0/I3742/net13	I0/I3742/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3744/T0	vdd	I0/I3744/net13	I0/I3744/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3733/T0	vdd	I0/I3733/net13	I0/I3733/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3747/T0	vdd	I0/I3747/net13	I0/I3747/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3741/T0	vdd	I0/I3741/net13	I0/I3741/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3745/T0	vdd	I0/I3745/net13	I0/I3745/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3758/T1	I0/I3758/net13	I0/I3758/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3759/T1	I0/I3759/net13	I0/I3759/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3766/T1	I0/I3766/net13	I0/I3766/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3768/T1	I0/I3768/net13	I0/I3768/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3774/T1	I0/I3774/net13	I0/I3774/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3776/T1	I0/I3776/net13	I0/I3776/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3765/T1	I0/I3765/net13	I0/I3765/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3779/T1	I0/I3779/net13	I0/I3779/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3773/T1	I0/I3773/net13	I0/I3773/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3777/T1	I0/I3777/net13	I0/I3777/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3758/T0	vdd	I0/I3758/net13	I0/I3758/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3759/T0	vdd	I0/I3759/net13	I0/I3759/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3766/T0	vdd	I0/I3766/net13	I0/I3766/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3768/T0	vdd	I0/I3768/net13	I0/I3768/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3774/T0	vdd	I0/I3774/net13	I0/I3774/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3776/T0	vdd	I0/I3776/net13	I0/I3776/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3765/T0	vdd	I0/I3765/net13	I0/I3765/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3779/T0	vdd	I0/I3779/net13	I0/I3779/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3773/T0	vdd	I0/I3773/net13	I0/I3773/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3777/T0	vdd	I0/I3777/net13	I0/I3777/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3534/T1	I0/I3534/net13	I0/I3534/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3535/T1	I0/I3535/net13	I0/I3535/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3542/T1	I0/I3542/net13	I0/I3542/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3544/T1	I0/I3544/net13	I0/I3544/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3550/T1	I0/I3550/net13	I0/I3550/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3552/T1	I0/I3552/net13	I0/I3552/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3541/T1	I0/I3541/net13	I0/I3541/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3555/T1	I0/I3555/net13	I0/I3555/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3549/T1	I0/I3549/net13	I0/I3549/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3553/T1	I0/I3553/net13	I0/I3553/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3534/T0	vdd	I0/I3534/net13	I0/I3534/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3535/T0	vdd	I0/I3535/net13	I0/I3535/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3542/T0	vdd	I0/I3542/net13	I0/I3542/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3544/T0	vdd	I0/I3544/net13	I0/I3544/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3550/T0	vdd	I0/I3550/net13	I0/I3550/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3552/T0	vdd	I0/I3552/net13	I0/I3552/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3541/T0	vdd	I0/I3541/net13	I0/I3541/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3555/T0	vdd	I0/I3555/net13	I0/I3555/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3549/T0	vdd	I0/I3549/net13	I0/I3549/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3553/T0	vdd	I0/I3553/net13	I0/I3553/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3566/T1	I0/I3566/net13	I0/I3566/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3567/T1	I0/I3567/net13	I0/I3567/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3574/T1	I0/I3574/net13	I0/I3574/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3576/T1	I0/I3576/net13	I0/I3576/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3582/T1	I0/I3582/net13	I0/I3582/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3584/T1	I0/I3584/net13	I0/I3584/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3573/T1	I0/I3573/net13	I0/I3573/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3587/T1	I0/I3587/net13	I0/I3587/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3581/T1	I0/I3581/net13	I0/I3581/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3585/T1	I0/I3585/net13	I0/I3585/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3566/T0	vdd	I0/I3566/net13	I0/I3566/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3567/T0	vdd	I0/I3567/net13	I0/I3567/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3574/T0	vdd	I0/I3574/net13	I0/I3574/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3576/T0	vdd	I0/I3576/net13	I0/I3576/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3582/T0	vdd	I0/I3582/net13	I0/I3582/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3584/T0	vdd	I0/I3584/net13	I0/I3584/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3573/T0	vdd	I0/I3573/net13	I0/I3573/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3587/T0	vdd	I0/I3587/net13	I0/I3587/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3581/T0	vdd	I0/I3581/net13	I0/I3581/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3585/T0	vdd	I0/I3585/net13	I0/I3585/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3598/T1	I0/I3598/net13	I0/I3598/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3599/T1	I0/I3599/net13	I0/I3599/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3606/T1	I0/I3606/net13	I0/I3606/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3608/T1	I0/I3608/net13	I0/I3608/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3614/T1	I0/I3614/net13	I0/I3614/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3616/T1	I0/I3616/net13	I0/I3616/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3605/T1	I0/I3605/net13	I0/I3605/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3619/T1	I0/I3619/net13	I0/I3619/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3613/T1	I0/I3613/net13	I0/I3613/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3617/T1	I0/I3617/net13	I0/I3617/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3598/T0	vdd	I0/I3598/net13	I0/I3598/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3599/T0	vdd	I0/I3599/net13	I0/I3599/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3606/T0	vdd	I0/I3606/net13	I0/I3606/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3608/T0	vdd	I0/I3608/net13	I0/I3608/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3614/T0	vdd	I0/I3614/net13	I0/I3614/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3616/T0	vdd	I0/I3616/net13	I0/I3616/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3605/T0	vdd	I0/I3605/net13	I0/I3605/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3619/T0	vdd	I0/I3619/net13	I0/I3619/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3613/T0	vdd	I0/I3613/net13	I0/I3613/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3617/T0	vdd	I0/I3617/net13	I0/I3617/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3630/T1	I0/I3630/net13	I0/I3630/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3631/T1	I0/I3631/net13	I0/I3631/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3638/T1	I0/I3638/net13	I0/I3638/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3640/T1	I0/I3640/net13	I0/I3640/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3646/T1	I0/I3646/net13	I0/I3646/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3648/T1	I0/I3648/net13	I0/I3648/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3637/T1	I0/I3637/net13	I0/I3637/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3651/T1	I0/I3651/net13	I0/I3651/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3645/T1	I0/I3645/net13	I0/I3645/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3649/T1	I0/I3649/net13	I0/I3649/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3630/T0	vdd	I0/I3630/net13	I0/I3630/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3631/T0	vdd	I0/I3631/net13	I0/I3631/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3638/T0	vdd	I0/I3638/net13	I0/I3638/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3640/T0	vdd	I0/I3640/net13	I0/I3640/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3646/T0	vdd	I0/I3646/net13	I0/I3646/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3648/T0	vdd	I0/I3648/net13	I0/I3648/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3637/T0	vdd	I0/I3637/net13	I0/I3637/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3651/T0	vdd	I0/I3651/net13	I0/I3651/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3645/T0	vdd	I0/I3645/net13	I0/I3645/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3649/T0	vdd	I0/I3649/net13	I0/I3649/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3406/T1	I0/I3406/net13	I0/I3406/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3407/T1	I0/I3407/net13	I0/I3407/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3414/T1	I0/I3414/net13	I0/I3414/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3416/T1	I0/I3416/net13	I0/I3416/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3422/T1	I0/I3422/net13	I0/I3422/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3424/T1	I0/I3424/net13	I0/I3424/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3413/T1	I0/I3413/net13	I0/I3413/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3427/T1	I0/I3427/net13	I0/I3427/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3421/T1	I0/I3421/net13	I0/I3421/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3425/T1	I0/I3425/net13	I0/I3425/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3406/T0	vdd	I0/I3406/net13	I0/I3406/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3407/T0	vdd	I0/I3407/net13	I0/I3407/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3414/T0	vdd	I0/I3414/net13	I0/I3414/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3416/T0	vdd	I0/I3416/net13	I0/I3416/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3422/T0	vdd	I0/I3422/net13	I0/I3422/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3424/T0	vdd	I0/I3424/net13	I0/I3424/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3413/T0	vdd	I0/I3413/net13	I0/I3413/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3427/T0	vdd	I0/I3427/net13	I0/I3427/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3421/T0	vdd	I0/I3421/net13	I0/I3421/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3425/T0	vdd	I0/I3425/net13	I0/I3425/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3757/T0	vdd	I0/I3757/net13	I0/I3757/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3743/T0	vdd	I0/I3743/net13	I0/I3743/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3754/T0	vdd	I0/I3754/net13	I0/I3754/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3753/T0	vdd	I0/I3753/net13	I0/I3753/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3757/T1	I0/I3757/net13	I0/I3757/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3743/T1	I0/I3743/net13	I0/I3743/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3754/T1	I0/I3754/net13	I0/I3754/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3753/T1	I0/I3753/net13	I0/I3753/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3789/T0	vdd	I0/I3789/net13	I0/I3789/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3775/T0	vdd	I0/I3775/net13	I0/I3775/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3786/T0	vdd	I0/I3786/net13	I0/I3786/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3785/T0	vdd	I0/I3785/net13	I0/I3785/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3789/T1	I0/I3789/net13	I0/I3789/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3775/T1	I0/I3775/net13	I0/I3775/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3786/T1	I0/I3786/net13	I0/I3786/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3785/T1	I0/I3785/net13	I0/I3785/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3565/T0	vdd	I0/I3565/net13	I0/I3565/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3551/T0	vdd	I0/I3551/net13	I0/I3551/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3562/T0	vdd	I0/I3562/net13	I0/I3562/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3561/T0	vdd	I0/I3561/net13	I0/I3561/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3565/T1	I0/I3565/net13	I0/I3565/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3551/T1	I0/I3551/net13	I0/I3551/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3562/T1	I0/I3562/net13	I0/I3562/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3561/T1	I0/I3561/net13	I0/I3561/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3597/T1	I0/I3597/net13	I0/I3597/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3583/T1	I0/I3583/net13	I0/I3583/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3594/T1	I0/I3594/net13	I0/I3594/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3593/T1	I0/I3593/net13	I0/I3593/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3597/T0	vdd	I0/I3597/net13	I0/I3597/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3583/T0	vdd	I0/I3583/net13	I0/I3583/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3594/T0	vdd	I0/I3594/net13	I0/I3594/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3593/T0	vdd	I0/I3593/net13	I0/I3593/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3629/T0	vdd	I0/I3629/net13	I0/I3629/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3615/T0	vdd	I0/I3615/net13	I0/I3615/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3626/T0	vdd	I0/I3626/net13	I0/I3626/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3625/T0	vdd	I0/I3625/net13	I0/I3625/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3629/T1	I0/I3629/net13	I0/I3629/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3615/T1	I0/I3615/net13	I0/I3615/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3626/T1	I0/I3626/net13	I0/I3626/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3625/T1	I0/I3625/net13	I0/I3625/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3661/T0	vdd	I0/I3661/net13	I0/I3661/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3647/T0	vdd	I0/I3647/net13	I0/I3647/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3658/T0	vdd	I0/I3658/net13	I0/I3658/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3657/T0	vdd	I0/I3657/net13	I0/I3657/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3661/T1	I0/I3661/net13	I0/I3661/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3647/T1	I0/I3647/net13	I0/I3647/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3658/T1	I0/I3658/net13	I0/I3658/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3657/T1	I0/I3657/net13	I0/I3657/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3437/T0	vdd	I0/I3437/net13	I0/I3437/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3423/T0	vdd	I0/I3423/net13	I0/I3423/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3434/T0	vdd	I0/I3434/net13	I0/I3434/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3433/T0	vdd	I0/I3433/net13	I0/I3433/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3437/T1	I0/I3437/net13	I0/I3437/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3423/T1	I0/I3423/net13	I0/I3423/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3434/T1	I0/I3434/net13	I0/I3434/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3433/T1	I0/I3433/net13	I0/I3433/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3570/T1	I0/I3570/net13	I0/I3570/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3538/T0	vdd	I0/I3538/net13	I0/I3538/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3538/T1	I0/I3538/net13	I0/I3538/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3762/T0	vdd	I0/I3762/net13	I0/I3762/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3762/T1	I0/I3762/net13	I0/I3762/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3730/T0	vdd	I0/I3730/net13	I0/I3730/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3730/T1	I0/I3730/net13	I0/I3730/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3410/T0	vdd	I0/I3410/net13	I0/I3410/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3410/T1	I0/I3410/net13	I0/I3410/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3634/T0	vdd	I0/I3634/net13	I0/I3634/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3634/T1	I0/I3634/net13	I0/I3634/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3602/T0	vdd	I0/I3602/net13	I0/I3602/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3602/T1	I0/I3602/net13	I0/I3602/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3570/T0	vdd	I0/I3570/net13	I0/I3570/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI80/T0	p6bar	y2bar	BL21bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI81/T0	BL21	y2bar	p6	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI82/T0	p6bar	y1bar	BL20bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI83/T0	BL20	y1bar	p6	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI84/T0	p7bar	y4bar	BL27bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI85/T0	BL27	y4bar	p7	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI86/T0	p7bar	y3bar	BL26bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI73/T0	BL17	y2bar	p5	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI74/T0	p5bar	y1bar	BL16bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI75/T0	BL16	y1bar	p5	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI76/T0	p6bar	y4bar	BL23bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI77/T0	BL23	y4bar	p6	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI78/T0	p6bar	y3bar	BL22bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI79/T0	BL22	y3bar	p6	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T0	vdd	I5/net24	I5/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T1	I5/net20	I5/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T9	vdd	I5/net20	I5/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI5/T10	data4	I5/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T10	I27/net23	data4	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T13	I27/net15	net681	p5	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T12	vdd	I27/net23	I27/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T14	I27/net7	p5	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI27/T15	p5bar	net681	I27/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T0	vdd	I6/net24	I6/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI6/T1	I6/net20	I6/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T1	I4/net20	I4/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T9	vdd	I4/net20	I4/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T10	data3	I4/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T10	I26/net23	data3	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T13	I26/net15	net681	p4	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T12	vdd	I26/net23	I26/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T14	I26/net7	p4	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI26/T15	p4bar	net681	I26/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI4/T0	vdd	I4/net24	I4/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI136/T1	vdd	clkout	BL17bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3452/T0	vdd	I0/I3452/net13	I0/I3452/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3444/T0	vdd	I0/I3444/net13	I0/I3444/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3443/T0	vdd	I0/I3443/net13	I0/I3443/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI136/T2	BL17	clkout	BL17bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI136/T0	BL17	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3452/T1	I0/I3452/net13	I0/I3452/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3444/T1	I0/I3444/net13	I0/I3444/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3443/T1	I0/I3443/net13	I0/I3443/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3468/T0	vdd	I0/I3468/net13	I0/I3468/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3449/T0	vdd	I0/I3449/net13	I0/I3449/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3464/T0	vdd	I0/I3464/net13	I0/I3464/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3462/T0	vdd	I0/I3462/net13	I0/I3462/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3468/T1	I0/I3468/net13	I0/I3468/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3449/T1	I0/I3449/net13	I0/I3449/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3464/T1	I0/I3464/net13	I0/I3464/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3462/T1	I0/I3462/net13	I0/I3462/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3458/T1	I0/I3458/net13	I0/I3458/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3450/T1	I0/I3450/net13	I0/I3450/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3451/T1	I0/I3451/net13	I0/I3451/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3441/T1	I0/I3441/net13	I0/I3441/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3467/T1	I0/I3467/net13	I0/I3467/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3461/T1	I0/I3461/net13	I0/I3461/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3447/T1	I0/I3447/net13	I0/I3447/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3440/T1	I0/I3440/net13	I0/I3440/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3463/T1	I0/I3463/net13	I0/I3463/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3460/T1	I0/I3460/net13	I0/I3460/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3458/T0	vdd	I0/I3458/net13	I0/I3458/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3450/T0	vdd	I0/I3450/net13	I0/I3450/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3451/T0	vdd	I0/I3451/net13	I0/I3451/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3441/T0	vdd	I0/I3441/net13	I0/I3441/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3467/T0	vdd	I0/I3467/net13	I0/I3467/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3461/T0	vdd	I0/I3461/net13	I0/I3461/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3447/T0	vdd	I0/I3447/net13	I0/I3447/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3440/T0	vdd	I0/I3440/net13	I0/I3440/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3463/T0	vdd	I0/I3463/net13	I0/I3463/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3460/T0	vdd	I0/I3460/net13	I0/I3460/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI137/T1	vdd	clkout	BL18bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3484/T0	vdd	I0/I3484/net13	I0/I3484/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3476/T0	vdd	I0/I3476/net13	I0/I3476/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3475/T0	vdd	I0/I3475/net13	I0/I3475/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI137/T2	BL18	clkout	BL18bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI137/T0	BL18	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3484/T1	I0/I3484/net13	I0/I3484/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3476/T1	I0/I3476/net13	I0/I3476/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3475/T1	I0/I3475/net13	I0/I3475/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3500/T0	vdd	I0/I3500/net13	I0/I3500/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3481/T0	vdd	I0/I3481/net13	I0/I3481/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3496/T0	vdd	I0/I3496/net13	I0/I3496/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3494/T0	vdd	I0/I3494/net13	I0/I3494/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3500/T1	I0/I3500/net13	I0/I3500/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3481/T1	I0/I3481/net13	I0/I3481/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3496/T1	I0/I3496/net13	I0/I3496/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3494/T1	I0/I3494/net13	I0/I3494/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3490/T1	I0/I3490/net13	I0/I3490/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3482/T1	I0/I3482/net13	I0/I3482/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3483/T1	I0/I3483/net13	I0/I3483/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3473/T1	I0/I3473/net13	I0/I3473/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3499/T1	I0/I3499/net13	I0/I3499/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3493/T1	I0/I3493/net13	I0/I3493/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3479/T1	I0/I3479/net13	I0/I3479/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3472/T1	I0/I3472/net13	I0/I3472/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3495/T1	I0/I3495/net13	I0/I3495/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3492/T1	I0/I3492/net13	I0/I3492/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3490/T0	vdd	I0/I3490/net13	I0/I3490/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3482/T0	vdd	I0/I3482/net13	I0/I3482/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3483/T0	vdd	I0/I3483/net13	I0/I3483/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3473/T0	vdd	I0/I3473/net13	I0/I3473/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3499/T0	vdd	I0/I3499/net13	I0/I3499/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3493/T0	vdd	I0/I3493/net13	I0/I3493/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3479/T0	vdd	I0/I3479/net13	I0/I3479/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3472/T0	vdd	I0/I3472/net13	I0/I3472/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3495/T0	vdd	I0/I3495/net13	I0/I3495/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3492/T0	vdd	I0/I3492/net13	I0/I3492/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI138/T1	vdd	clkout	BL19bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3516/T0	vdd	I0/I3516/net13	I0/I3516/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3508/T0	vdd	I0/I3508/net13	I0/I3508/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3507/T0	vdd	I0/I3507/net13	I0/I3507/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI138/T2	BL19	clkout	BL19bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI138/T0	BL19	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3516/T1	I0/I3516/net13	I0/I3516/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3508/T1	I0/I3508/net13	I0/I3508/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3507/T1	I0/I3507/net13	I0/I3507/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3532/T0	vdd	I0/I3532/net13	I0/I3532/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3513/T0	vdd	I0/I3513/net13	I0/I3513/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3528/T0	vdd	I0/I3528/net13	I0/I3528/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3526/T0	vdd	I0/I3526/net13	I0/I3526/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3532/T1	I0/I3532/net13	I0/I3532/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3513/T1	I0/I3513/net13	I0/I3513/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3528/T1	I0/I3528/net13	I0/I3528/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3526/T1	I0/I3526/net13	I0/I3526/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3522/T1	I0/I3522/net13	I0/I3522/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3514/T1	I0/I3514/net13	I0/I3514/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3515/T1	I0/I3515/net13	I0/I3515/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3505/T1	I0/I3505/net13	I0/I3505/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3531/T1	I0/I3531/net13	I0/I3531/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3525/T1	I0/I3525/net13	I0/I3525/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3511/T1	I0/I3511/net13	I0/I3511/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3504/T1	I0/I3504/net13	I0/I3504/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3527/T1	I0/I3527/net13	I0/I3527/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3524/T1	I0/I3524/net13	I0/I3524/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3522/T0	vdd	I0/I3522/net13	I0/I3522/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3514/T0	vdd	I0/I3514/net13	I0/I3514/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3515/T0	vdd	I0/I3515/net13	I0/I3515/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3505/T0	vdd	I0/I3505/net13	I0/I3505/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3531/T0	vdd	I0/I3531/net13	I0/I3531/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3525/T0	vdd	I0/I3525/net13	I0/I3525/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3511/T0	vdd	I0/I3511/net13	I0/I3511/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3504/T0	vdd	I0/I3504/net13	I0/I3504/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3527/T0	vdd	I0/I3527/net13	I0/I3527/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3524/T0	vdd	I0/I3524/net13	I0/I3524/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI131/T1	vdd	clkout	BL12bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3292/T0	vdd	I0/I3292/net13	I0/I3292/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3284/T0	vdd	I0/I3284/net13	I0/I3284/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3283/T0	vdd	I0/I3283/net13	I0/I3283/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI131/T2	BL12	clkout	BL12bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI131/T0	BL12	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3292/T1	I0/I3292/net13	I0/I3292/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3284/T1	I0/I3284/net13	I0/I3284/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3283/T1	I0/I3283/net13	I0/I3283/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3308/T0	vdd	I0/I3308/net13	I0/I3308/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3289/T0	vdd	I0/I3289/net13	I0/I3289/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3304/T0	vdd	I0/I3304/net13	I0/I3304/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3302/T0	vdd	I0/I3302/net13	I0/I3302/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3308/T1	I0/I3308/net13	I0/I3308/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3289/T1	I0/I3289/net13	I0/I3289/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3304/T1	I0/I3304/net13	I0/I3304/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3302/T1	I0/I3302/net13	I0/I3302/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3298/T1	I0/I3298/net13	I0/I3298/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3290/T1	I0/I3290/net13	I0/I3290/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3291/T1	I0/I3291/net13	I0/I3291/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3281/T1	I0/I3281/net13	I0/I3281/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3307/T1	I0/I3307/net13	I0/I3307/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3301/T1	I0/I3301/net13	I0/I3301/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3287/T1	I0/I3287/net13	I0/I3287/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3280/T1	I0/I3280/net13	I0/I3280/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3303/T1	I0/I3303/net13	I0/I3303/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3300/T1	I0/I3300/net13	I0/I3300/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3298/T0	vdd	I0/I3298/net13	I0/I3298/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3290/T0	vdd	I0/I3290/net13	I0/I3290/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3291/T0	vdd	I0/I3291/net13	I0/I3291/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3281/T0	vdd	I0/I3281/net13	I0/I3281/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3307/T0	vdd	I0/I3307/net13	I0/I3307/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3301/T0	vdd	I0/I3301/net13	I0/I3301/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3287/T0	vdd	I0/I3287/net13	I0/I3287/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3280/T0	vdd	I0/I3280/net13	I0/I3280/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3303/T0	vdd	I0/I3303/net13	I0/I3303/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3300/T0	vdd	I0/I3300/net13	I0/I3300/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3438/T1	I0/I3438/net13	I0/I3438/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3439/T1	I0/I3439/net13	I0/I3439/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3446/T1	I0/I3446/net13	I0/I3446/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3448/T1	I0/I3448/net13	I0/I3448/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3454/T1	I0/I3454/net13	I0/I3454/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3456/T1	I0/I3456/net13	I0/I3456/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3445/T1	I0/I3445/net13	I0/I3445/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3459/T1	I0/I3459/net13	I0/I3459/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3453/T1	I0/I3453/net13	I0/I3453/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3457/T1	I0/I3457/net13	I0/I3457/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3438/T0	vdd	I0/I3438/net13	I0/I3438/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3439/T0	vdd	I0/I3439/net13	I0/I3439/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3446/T0	vdd	I0/I3446/net13	I0/I3446/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3448/T0	vdd	I0/I3448/net13	I0/I3448/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3454/T0	vdd	I0/I3454/net13	I0/I3454/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3456/T0	vdd	I0/I3456/net13	I0/I3456/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3445/T0	vdd	I0/I3445/net13	I0/I3445/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3459/T0	vdd	I0/I3459/net13	I0/I3459/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3453/T0	vdd	I0/I3453/net13	I0/I3453/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3457/T0	vdd	I0/I3457/net13	I0/I3457/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3470/T1	I0/I3470/net13	I0/I3470/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3471/T1	I0/I3471/net13	I0/I3471/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3478/T1	I0/I3478/net13	I0/I3478/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3480/T1	I0/I3480/net13	I0/I3480/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3486/T1	I0/I3486/net13	I0/I3486/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3488/T1	I0/I3488/net13	I0/I3488/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3477/T1	I0/I3477/net13	I0/I3477/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3491/T1	I0/I3491/net13	I0/I3491/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3485/T1	I0/I3485/net13	I0/I3485/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3489/T1	I0/I3489/net13	I0/I3489/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3470/T0	vdd	I0/I3470/net13	I0/I3470/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3471/T0	vdd	I0/I3471/net13	I0/I3471/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3478/T0	vdd	I0/I3478/net13	I0/I3478/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3480/T0	vdd	I0/I3480/net13	I0/I3480/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3486/T0	vdd	I0/I3486/net13	I0/I3486/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3488/T0	vdd	I0/I3488/net13	I0/I3488/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3477/T0	vdd	I0/I3477/net13	I0/I3477/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3491/T0	vdd	I0/I3491/net13	I0/I3491/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3485/T0	vdd	I0/I3485/net13	I0/I3485/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3489/T0	vdd	I0/I3489/net13	I0/I3489/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3502/T1	I0/I3502/net13	I0/I3502/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3503/T1	I0/I3503/net13	I0/I3503/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3510/T1	I0/I3510/net13	I0/I3510/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3512/T1	I0/I3512/net13	I0/I3512/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3518/T1	I0/I3518/net13	I0/I3518/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3520/T1	I0/I3520/net13	I0/I3520/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3509/T1	I0/I3509/net13	I0/I3509/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3523/T1	I0/I3523/net13	I0/I3523/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3517/T1	I0/I3517/net13	I0/I3517/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3521/T1	I0/I3521/net13	I0/I3521/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3502/T0	vdd	I0/I3502/net13	I0/I3502/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3503/T0	vdd	I0/I3503/net13	I0/I3503/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3510/T0	vdd	I0/I3510/net13	I0/I3510/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3512/T0	vdd	I0/I3512/net13	I0/I3512/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3518/T0	vdd	I0/I3518/net13	I0/I3518/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3520/T0	vdd	I0/I3520/net13	I0/I3520/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3509/T0	vdd	I0/I3509/net13	I0/I3509/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3523/T0	vdd	I0/I3523/net13	I0/I3523/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3517/T0	vdd	I0/I3517/net13	I0/I3517/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3521/T0	vdd	I0/I3521/net13	I0/I3521/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3278/T1	I0/I3278/net13	I0/I3278/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3279/T1	I0/I3279/net13	I0/I3279/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3286/T1	I0/I3286/net13	I0/I3286/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3288/T1	I0/I3288/net13	I0/I3288/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3294/T1	I0/I3294/net13	I0/I3294/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3296/T1	I0/I3296/net13	I0/I3296/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3285/T1	I0/I3285/net13	I0/I3285/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3299/T1	I0/I3299/net13	I0/I3299/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3293/T1	I0/I3293/net13	I0/I3293/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3297/T1	I0/I3297/net13	I0/I3297/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3278/T0	vdd	I0/I3278/net13	I0/I3278/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3279/T0	vdd	I0/I3279/net13	I0/I3279/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3286/T0	vdd	I0/I3286/net13	I0/I3286/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3288/T0	vdd	I0/I3288/net13	I0/I3288/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3294/T0	vdd	I0/I3294/net13	I0/I3294/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3296/T0	vdd	I0/I3296/net13	I0/I3296/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3285/T0	vdd	I0/I3285/net13	I0/I3285/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3299/T0	vdd	I0/I3299/net13	I0/I3299/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3293/T0	vdd	I0/I3293/net13	I0/I3293/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3297/T0	vdd	I0/I3297/net13	I0/I3297/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3469/T0	vdd	I0/I3469/net13	I0/I3469/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3455/T0	vdd	I0/I3455/net13	I0/I3455/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3466/T0	vdd	I0/I3466/net13	I0/I3466/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3465/T0	vdd	I0/I3465/net13	I0/I3465/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3442/T0	vdd	I0/I3442/net13	I0/I3442/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3469/T1	I0/I3469/net13	I0/I3469/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3455/T1	I0/I3455/net13	I0/I3455/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3466/T1	I0/I3466/net13	I0/I3466/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3465/T1	I0/I3465/net13	I0/I3465/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3442/T1	I0/I3442/net13	I0/I3442/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3501/T0	vdd	I0/I3501/net13	I0/I3501/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3487/T0	vdd	I0/I3487/net13	I0/I3487/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3498/T0	vdd	I0/I3498/net13	I0/I3498/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3497/T0	vdd	I0/I3497/net13	I0/I3497/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3474/T0	vdd	I0/I3474/net13	I0/I3474/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3501/T1	I0/I3501/net13	I0/I3501/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3487/T1	I0/I3487/net13	I0/I3487/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3498/T1	I0/I3498/net13	I0/I3498/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3497/T1	I0/I3497/net13	I0/I3497/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3474/T1	I0/I3474/net13	I0/I3474/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3533/T0	vdd	I0/I3533/net13	I0/I3533/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3519/T0	vdd	I0/I3519/net13	I0/I3519/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3530/T0	vdd	I0/I3530/net13	I0/I3530/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3529/T0	vdd	I0/I3529/net13	I0/I3529/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3506/T0	vdd	I0/I3506/net13	I0/I3506/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3533/T1	I0/I3533/net13	I0/I3533/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3519/T1	I0/I3519/net13	I0/I3519/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3530/T1	I0/I3530/net13	I0/I3530/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3529/T1	I0/I3529/net13	I0/I3529/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3506/T1	I0/I3506/net13	I0/I3506/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3309/T0	vdd	I0/I3309/net13	I0/I3309/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3295/T0	vdd	I0/I3295/net13	I0/I3295/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3306/T0	vdd	I0/I3306/net13	I0/I3306/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3305/T0	vdd	I0/I3305/net13	I0/I3305/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3282/T0	vdd	I0/I3282/net13	I0/I3282/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3309/T1	I0/I3309/net13	I0/I3309/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3295/T1	I0/I3295/net13	I0/I3295/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3306/T1	I0/I3306/net13	I0/I3306/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3305/T1	I0/I3305/net13	I0/I3305/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3282/T1	I0/I3282/net13	I0/I3282/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI67/T0	BL12	y1bar	p4	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI68/T0	p5bar	y4bar	BL19bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI69/T0	BL19	y4bar	p5	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI70/T0	p5bar	y3bar	BL18bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI71/T0	BL18	y3bar	p5	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI72/T0	p5bar	y2bar	BL17bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T9	vdd	I3/net20	I3/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T10	data2	I3/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T10	I25/net23	data2	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T13	I25/net15	net681	net740	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T12	vdd	I25/net23	I25/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=7.2e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T14	I25/net7	net740	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=7.2e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI25/T15	net741	net681	I25/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=7.2e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T17	I30/net57	I30/net61	vdd	vdd	pfet	L=0.12U
+ W=2.44U
+ AD=0.7808P	AS=0.7808P	PD=5.52U	PS=5.52U
+ wt=2.44e-06 wf=2.44e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=3.288e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.68e-14 nrs=0.091858 nrd=0.091858 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI66/T0	p4bar	y1bar	BL12bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T18	net681	I30/net57	vdd	vdd	pfet	L=0.12U
+ W=9U
+ AD=2.88P	AS=2.88P	PD=18.64U	PS=18.64U
+ wt=9e-06 wf=9e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.104e-12 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0245673 nrd=0.0245673 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI133/T0	BL14	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3356/T1	I0/I3356/net13	I0/I3356/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI132/T1	vdd	clkout	BL13bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3324/T0	vdd	I0/I3324/net13	I0/I3324/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI132/T2	BL13	clkout	BL13bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI132/T0	BL13	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3324/T1	I0/I3324/net13	I0/I3324/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI133/T2	BL14	clkout	BL14bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI134/T1	vdd	clkout	BL15bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3388/T0	vdd	I0/I3388/net13	I0/I3388/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI134/T2	BL15	clkout	BL15bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI134/T0	BL15	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3388/T1	I0/I3388/net13	I0/I3388/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI133/T1	vdd	clkout	BL14bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3356/T0	vdd	I0/I3356/net13	I0/I3356/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3348/T1	I0/I3348/net13	I0/I3348/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3347/T1	I0/I3347/net13	I0/I3347/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3316/T0	vdd	I0/I3316/net13	I0/I3316/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3315/T0	vdd	I0/I3315/net13	I0/I3315/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3316/T1	I0/I3316/net13	I0/I3316/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3315/T1	I0/I3315/net13	I0/I3315/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3380/T0	vdd	I0/I3380/net13	I0/I3380/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3379/T0	vdd	I0/I3379/net13	I0/I3379/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3380/T1	I0/I3380/net13	I0/I3380/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3379/T1	I0/I3379/net13	I0/I3379/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3348/T0	vdd	I0/I3348/net13	I0/I3348/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3347/T0	vdd	I0/I3347/net13	I0/I3347/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3340/T0	vdd	I0/I3340/net13	I0/I3340/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3321/T0	vdd	I0/I3321/net13	I0/I3321/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3336/T0	vdd	I0/I3336/net13	I0/I3336/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3334/T0	vdd	I0/I3334/net13	I0/I3334/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3340/T1	I0/I3340/net13	I0/I3340/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3321/T1	I0/I3321/net13	I0/I3321/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3336/T1	I0/I3336/net13	I0/I3336/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3334/T1	I0/I3334/net13	I0/I3334/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3372/T1	I0/I3372/net13	I0/I3372/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3353/T1	I0/I3353/net13	I0/I3353/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3368/T1	I0/I3368/net13	I0/I3368/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3366/T1	I0/I3366/net13	I0/I3366/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3372/T0	vdd	I0/I3372/net13	I0/I3372/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3353/T0	vdd	I0/I3353/net13	I0/I3353/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3368/T0	vdd	I0/I3368/net13	I0/I3368/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3366/T0	vdd	I0/I3366/net13	I0/I3366/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3404/T0	vdd	I0/I3404/net13	I0/I3404/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3385/T0	vdd	I0/I3385/net13	I0/I3385/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3400/T0	vdd	I0/I3400/net13	I0/I3400/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3398/T0	vdd	I0/I3398/net13	I0/I3398/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3404/T1	I0/I3404/net13	I0/I3404/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3385/T1	I0/I3385/net13	I0/I3385/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3400/T1	I0/I3400/net13	I0/I3400/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3398/T1	I0/I3398/net13	I0/I3398/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3330/T1	I0/I3330/net13	I0/I3330/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3322/T1	I0/I3322/net13	I0/I3322/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3323/T1	I0/I3323/net13	I0/I3323/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3313/T1	I0/I3313/net13	I0/I3313/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3339/T1	I0/I3339/net13	I0/I3339/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3333/T1	I0/I3333/net13	I0/I3333/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3319/T1	I0/I3319/net13	I0/I3319/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3312/T1	I0/I3312/net13	I0/I3312/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3335/T1	I0/I3335/net13	I0/I3335/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3332/T1	I0/I3332/net13	I0/I3332/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3330/T0	vdd	I0/I3330/net13	I0/I3330/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3322/T0	vdd	I0/I3322/net13	I0/I3322/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3323/T0	vdd	I0/I3323/net13	I0/I3323/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3313/T0	vdd	I0/I3313/net13	I0/I3313/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3339/T0	vdd	I0/I3339/net13	I0/I3339/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3333/T0	vdd	I0/I3333/net13	I0/I3333/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3319/T0	vdd	I0/I3319/net13	I0/I3319/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3312/T0	vdd	I0/I3312/net13	I0/I3312/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3335/T0	vdd	I0/I3335/net13	I0/I3335/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3332/T0	vdd	I0/I3332/net13	I0/I3332/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3362/T1	I0/I3362/net13	I0/I3362/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3354/T1	I0/I3354/net13	I0/I3354/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3355/T1	I0/I3355/net13	I0/I3355/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3345/T1	I0/I3345/net13	I0/I3345/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3371/T1	I0/I3371/net13	I0/I3371/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3365/T1	I0/I3365/net13	I0/I3365/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3351/T1	I0/I3351/net13	I0/I3351/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3344/T1	I0/I3344/net13	I0/I3344/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3367/T1	I0/I3367/net13	I0/I3367/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3364/T1	I0/I3364/net13	I0/I3364/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3362/T0	vdd	I0/I3362/net13	I0/I3362/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3354/T0	vdd	I0/I3354/net13	I0/I3354/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3355/T0	vdd	I0/I3355/net13	I0/I3355/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3345/T0	vdd	I0/I3345/net13	I0/I3345/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3371/T0	vdd	I0/I3371/net13	I0/I3371/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3365/T0	vdd	I0/I3365/net13	I0/I3365/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3351/T0	vdd	I0/I3351/net13	I0/I3351/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3344/T0	vdd	I0/I3344/net13	I0/I3344/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3367/T0	vdd	I0/I3367/net13	I0/I3367/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3364/T0	vdd	I0/I3364/net13	I0/I3364/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3394/T1	I0/I3394/net13	I0/I3394/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3386/T1	I0/I3386/net13	I0/I3386/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3387/T1	I0/I3387/net13	I0/I3387/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3377/T1	I0/I3377/net13	I0/I3377/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3403/T1	I0/I3403/net13	I0/I3403/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3397/T1	I0/I3397/net13	I0/I3397/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3383/T1	I0/I3383/net13	I0/I3383/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3376/T1	I0/I3376/net13	I0/I3376/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3399/T1	I0/I3399/net13	I0/I3399/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3396/T1	I0/I3396/net13	I0/I3396/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3394/T0	vdd	I0/I3394/net13	I0/I3394/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3386/T0	vdd	I0/I3386/net13	I0/I3386/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3387/T0	vdd	I0/I3387/net13	I0/I3387/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3377/T0	vdd	I0/I3377/net13	I0/I3377/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3403/T0	vdd	I0/I3403/net13	I0/I3403/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3397/T0	vdd	I0/I3397/net13	I0/I3397/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3383/T0	vdd	I0/I3383/net13	I0/I3383/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3376/T0	vdd	I0/I3376/net13	I0/I3376/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3399/T0	vdd	I0/I3399/net13	I0/I3399/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3396/T0	vdd	I0/I3396/net13	I0/I3396/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3310/T1	I0/I3310/net13	I0/I3310/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3311/T1	I0/I3311/net13	I0/I3311/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3318/T1	I0/I3318/net13	I0/I3318/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3320/T1	I0/I3320/net13	I0/I3320/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3326/T1	I0/I3326/net13	I0/I3326/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3328/T1	I0/I3328/net13	I0/I3328/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3317/T1	I0/I3317/net13	I0/I3317/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3331/T1	I0/I3331/net13	I0/I3331/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3325/T1	I0/I3325/net13	I0/I3325/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3329/T1	I0/I3329/net13	I0/I3329/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3310/T0	vdd	I0/I3310/net13	I0/I3310/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3311/T0	vdd	I0/I3311/net13	I0/I3311/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3318/T0	vdd	I0/I3318/net13	I0/I3318/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3320/T0	vdd	I0/I3320/net13	I0/I3320/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3326/T0	vdd	I0/I3326/net13	I0/I3326/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3328/T0	vdd	I0/I3328/net13	I0/I3328/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3317/T0	vdd	I0/I3317/net13	I0/I3317/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3331/T0	vdd	I0/I3331/net13	I0/I3331/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3325/T0	vdd	I0/I3325/net13	I0/I3325/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3329/T0	vdd	I0/I3329/net13	I0/I3329/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3342/T1	I0/I3342/net13	I0/I3342/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3343/T1	I0/I3343/net13	I0/I3343/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3350/T1	I0/I3350/net13	I0/I3350/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3352/T1	I0/I3352/net13	I0/I3352/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3358/T1	I0/I3358/net13	I0/I3358/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3360/T1	I0/I3360/net13	I0/I3360/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3349/T1	I0/I3349/net13	I0/I3349/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3363/T1	I0/I3363/net13	I0/I3363/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3357/T1	I0/I3357/net13	I0/I3357/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3361/T1	I0/I3361/net13	I0/I3361/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3342/T0	vdd	I0/I3342/net13	I0/I3342/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3343/T0	vdd	I0/I3343/net13	I0/I3343/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3350/T0	vdd	I0/I3350/net13	I0/I3350/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3352/T0	vdd	I0/I3352/net13	I0/I3352/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3358/T0	vdd	I0/I3358/net13	I0/I3358/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3360/T0	vdd	I0/I3360/net13	I0/I3360/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3349/T0	vdd	I0/I3349/net13	I0/I3349/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3363/T0	vdd	I0/I3363/net13	I0/I3363/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3357/T0	vdd	I0/I3357/net13	I0/I3357/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3361/T0	vdd	I0/I3361/net13	I0/I3361/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3374/T1	I0/I3374/net13	I0/I3374/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3375/T1	I0/I3375/net13	I0/I3375/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3382/T1	I0/I3382/net13	I0/I3382/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3384/T1	I0/I3384/net13	I0/I3384/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3390/T1	I0/I3390/net13	I0/I3390/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3392/T1	I0/I3392/net13	I0/I3392/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3381/T1	I0/I3381/net13	I0/I3381/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3395/T1	I0/I3395/net13	I0/I3395/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3389/T1	I0/I3389/net13	I0/I3389/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3393/T1	I0/I3393/net13	I0/I3393/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3374/T0	vdd	I0/I3374/net13	I0/I3374/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3375/T0	vdd	I0/I3375/net13	I0/I3375/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3382/T0	vdd	I0/I3382/net13	I0/I3382/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3384/T0	vdd	I0/I3384/net13	I0/I3384/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3390/T0	vdd	I0/I3390/net13	I0/I3390/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3392/T0	vdd	I0/I3392/net13	I0/I3392/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3381/T0	vdd	I0/I3381/net13	I0/I3381/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3395/T0	vdd	I0/I3395/net13	I0/I3395/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3389/T0	vdd	I0/I3389/net13	I0/I3389/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3393/T0	vdd	I0/I3393/net13	I0/I3393/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3341/T0	vdd	I0/I3341/net13	I0/I3341/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3327/T0	vdd	I0/I3327/net13	I0/I3327/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3338/T0	vdd	I0/I3338/net13	I0/I3338/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3337/T0	vdd	I0/I3337/net13	I0/I3337/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3314/T0	vdd	I0/I3314/net13	I0/I3314/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3341/T1	I0/I3341/net13	I0/I3341/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3327/T1	I0/I3327/net13	I0/I3327/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3338/T1	I0/I3338/net13	I0/I3338/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3337/T1	I0/I3337/net13	I0/I3337/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3314/T1	I0/I3314/net13	I0/I3314/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3373/T1	I0/I3373/net13	I0/I3373/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3359/T1	I0/I3359/net13	I0/I3359/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3370/T1	I0/I3370/net13	I0/I3370/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3369/T1	I0/I3369/net13	I0/I3369/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3346/T1	I0/I3346/net13	I0/I3346/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3373/T0	vdd	I0/I3373/net13	I0/I3373/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3359/T0	vdd	I0/I3359/net13	I0/I3359/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3370/T0	vdd	I0/I3370/net13	I0/I3370/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3369/T0	vdd	I0/I3369/net13	I0/I3369/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3346/T0	vdd	I0/I3346/net13	I0/I3346/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3405/T0	vdd	I0/I3405/net13	I0/I3405/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3391/T0	vdd	I0/I3391/net13	I0/I3391/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3402/T0	vdd	I0/I3402/net13	I0/I3402/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3401/T0	vdd	I0/I3401/net13	I0/I3401/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3378/T0	vdd	I0/I3378/net13	I0/I3378/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3405/T1	I0/I3405/net13	I0/I3405/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3391/T1	I0/I3391/net13	I0/I3391/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3402/T1	I0/I3402/net13	I0/I3402/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3401/T1	I0/I3401/net13	I0/I3401/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3378/T1	I0/I3378/net13	I0/I3378/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI59/T0	BL8	y1bar	net740	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI60/T0	p4bar	y4bar	BL15bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI61/T0	BL15	y4bar	p4	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI62/T0	p4bar	y3bar	BL14bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI63/T0	BL14	y3bar	p4	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI64/T0	p4bar	y2bar	BL13bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI65/T0	BL13	y2bar	p4	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T14	I24/net7	net262	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T15	net256	net681	I24/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T10	I30/net49	wr	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.32e-14 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI3/T0	vdd	I3/net24	I3/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI3/T1	I3/net20	I3/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T7	I30/net61	wr	vdd	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.32e-14 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI2/T9	vdd	I2/net20	I2/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T10	data1	I2/net8	vdd	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T23	I30/net17	I30/net49	vdd	vdd	pfet	L=0.12U
+ W=1.28U
+ AD=0.4096P	AS=0.4096P	PD=3.2U	PS=3.2U
+ wt=1.28e-06 wf=1.28e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=4.72e-14 nrs=0.178138 nrd=0.178138 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI24/T10	I24/net23	data1	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T13	I24/net15	net681	net262	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI24/T12	vdd	I24/net23	I24/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T25	net680	I30/net41	vdd	vdd	pfet	L=0.12U
+ W=9U
+ AD=2.88P	AS=2.88P	PD=18.64U	PS=18.64U
+ wt=9e-06 wf=9e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.104e-12 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=4.8e-15 panw10=7.2e-14 nrs=0.0245673 nrd=0.0245673 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI128/T0	BL9	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3132/T1	I0/I3132/net13	I0/I3132/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI127/T1	vdd	clkout	BL8bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3100/T0	vdd	I0/I3100/net13	I0/I3100/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI127/T2	BL8	clkout	BL8bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI127/T0	BL8	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3100/T1	I0/I3100/net13	I0/I3100/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI128/T2	BL9	clkout	BL9bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI129/T1	vdd	clkout	BL10bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3164/T0	vdd	I0/I3164/net13	I0/I3164/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI129/T2	BL10	clkout	BL10bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI129/T0	BL10	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3164/T1	I0/I3164/net13	I0/I3164/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI128/T1	vdd	clkout	BL9bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3132/T0	vdd	I0/I3132/net13	I0/I3132/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3124/T1	I0/I3124/net13	I0/I3124/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3123/T1	I0/I3123/net13	I0/I3123/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3092/T0	vdd	I0/I3092/net13	I0/I3092/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3091/T0	vdd	I0/I3091/net13	I0/I3091/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3092/T1	I0/I3092/net13	I0/I3092/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3091/T1	I0/I3091/net13	I0/I3091/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3156/T0	vdd	I0/I3156/net13	I0/I3156/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3155/T0	vdd	I0/I3155/net13	I0/I3155/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3156/T1	I0/I3156/net13	I0/I3156/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3155/T1	I0/I3155/net13	I0/I3155/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3124/T0	vdd	I0/I3124/net13	I0/I3124/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3123/T0	vdd	I0/I3123/net13	I0/I3123/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI123/T0	BL4	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I107/T1	I0/I107/net13	I0/I107/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI130/T1	vdd	clkout	BL11bar	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3196/T0	vdd	I0/I3196/net13	I0/I3196/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI130/T2	BL11	clkout	BL11bar	vdd	pfet	L=0.12U
+ W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI130/T0	BL11	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3196/T1	I0/I3196/net13	I0/I3196/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI123/T2	BL4	clkout	BL4bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI124/T1	vdd	clkout	BL5bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3004/T0	vdd	I0/I3004/net13	I0/I3004/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI124/T2	BL5	clkout	BL5bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI124/T0	BL5	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3004/T1	I0/I3004/net13	I0/I3004/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI123/T1	vdd	clkout	BL4bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I107/T0	vdd	I0/I107/net13	I0/I107/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I115/T1	I0/I115/net13	I0/I115/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I116/T1	I0/I116/net13	I0/I116/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3188/T0	vdd	I0/I3188/net13	I0/I3188/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3187/T0	vdd	I0/I3187/net13	I0/I3187/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3188/T1	I0/I3188/net13	I0/I3188/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3187/T1	I0/I3187/net13	I0/I3187/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2996/T0	vdd	I0/I2996/net13	I0/I2996/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2995/T0	vdd	I0/I2995/net13	I0/I2995/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2996/T1	I0/I2996/net13	I0/I2996/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2995/T1	I0/I2995/net13	I0/I2995/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I115/T0	vdd	I0/I115/net13	I0/I115/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I116/T0	vdd	I0/I116/net13	I0/I116/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI126/T0	BL7	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3068/T1	I0/I3068/net13	I0/I3068/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI125/T1	vdd	clkout	BL6bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3036/T0	vdd	I0/I3036/net13	I0/I3036/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI125/T2	BL6	clkout	BL6bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI125/T0	BL6	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3036/T1	I0/I3036/net13	I0/I3036/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI126/T2	BL7	clkout	BL7bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI119/T1	vdd	clkout	BL0bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I84/T0	vdd	I0/I84/net13	I0/I84/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI119/T2	BL0	clkout	BL0bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI119/T0	BL0	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I84/T1	I0/I84/net13	I0/I84/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI126/T1	vdd	clkout	BL7bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3068/T0	vdd	I0/I3068/net13	I0/I3068/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3060/T1	I0/I3060/net13	I0/I3060/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3059/T1	I0/I3059/net13	I0/I3059/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3028/T0	vdd	I0/I3028/net13	I0/I3028/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3027/T0	vdd	I0/I3027/net13	I0/I3027/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3028/T1	I0/I3028/net13	I0/I3028/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3027/T1	I0/I3027/net13	I0/I3027/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I82/T0	vdd	I0/I82/net13	I0/I82/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I6/T0	vdd	I0/I6/net13	I0/I6/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I82/T1	I0/I82/net13	I0/I82/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I6/T1	I0/I6/net13	I0/I6/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3060/T0	vdd	I0/I3060/net13	I0/I3060/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3059/T0	vdd	I0/I3059/net13	I0/I3059/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI121/T0	BL2	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2894/T1	I0/I2894/net13	I0/I2894/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI120/T1	vdd	clkout	BL1bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2862/T0	vdd	I0/I2862/net13	I0/I2862/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI120/T2	BL1	clkout	BL1bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI120/T0	BL1	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2862/T1	I0/I2862/net13	I0/I2862/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI121/T2	BL2	clkout	BL2bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI122/T1	vdd	clkout	BL3bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw8=7.68e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2926/T0	vdd	I0/I2926/net13	I0/I2926/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI122/T2	BL3	clkout	BL3bar	vdd	pfet	L=0.12U	W=0.6U
+ AD=0.342P	AS=0.33P	PD=2.34U	PS=2.3U
+ wt=6e-07 wf=6e-07 sd=0 sb=5.7e-07 sa=5.5e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=7.2e-14 panw8=1.2e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.396396 nrd=0.396396 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI122/T0	BL3	clkout	vdd	vdd	pfet	L=0.12U	W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=7.76e-14 panw10=1.312e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2926/T1	I0/I2926/net13	I0/I2926/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI121/T1	vdd	clkout	BL2bar	vdd	pfet	L=0.12U	W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.64e-14 panw10=1.056e-13 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2894/T0	vdd	I0/I2894/net13	I0/I2894/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2895/T1	I0/I2895/net13	I0/I2895/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2909/T1	I0/I2909/net13	I0/I2909/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2866/T0	vdd	I0/I2866/net13	I0/I2866/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2888/T0	vdd	I0/I2888/net13	I0/I2888/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2866/T1	I0/I2866/net13	I0/I2866/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2888/T1	I0/I2888/net13	I0/I2888/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2934/T0	vdd	I0/I2934/net13	I0/I2934/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2933/T0	vdd	I0/I2933/net13	I0/I2933/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2934/T1	I0/I2934/net13	I0/I2934/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.4e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.96e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2933/T1	I0/I2933/net13	I0/I2933/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.4e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.96e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2895/T0	vdd	I0/I2895/net13	I0/I2895/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2909/T0	vdd	I0/I2909/net13	I0/I2909/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI159/T3	vdd	I159/net28	clkout	vdd	pfet	L=0.12U
+ W=34.58U
+ AD=11.0656P	AS=11.0656P	PD=69.8U	PS=69.8U
+ wt=3.458e-05 wf=3.458e-05 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=3.8112e-12 panw10=5.88e-14 nrs=0.00637035 nrd=0.00637035 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T5	vdd	I1/net176	I1/net1308	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T4	I1/net1308	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T76	vdd	I1/net112	I1/net1260	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T75	I1/net1260	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T79	vdd	I1/net76	I1/net1220	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T80	I1/net1220	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T0	net955	I1/net1308	vdd	vdd	pfet	L=0.12U	W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T77	net954	I1/net1260	vdd	vdd	pfet	L=0.12U	W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T78	net953	I1/net1220	vdd	vdd	pfet	L=0.12U	W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T6	I1/net176	I1/net1292	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T74	I1/net112	I1/net1248	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T81	I1/net76	I1/net1208	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T13	vdd	I1/net160	I1/net1292	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T12	I1/net1292	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T11	vdd	I1/a4bar	I1/net1292	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T73	vdd	I1/net160	I1/net1248	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T72	I1/net1248	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T71	vdd	I1/a4	I1/net1248	vdd	pfet	L=0.12U	W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T82	vdd	I1/net160	I1/net1208	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T83	I1/net1208	I1/a3	vdd	vdd	pfet	L=0.12U	W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T84	vdd	I1/a4bar	I1/net1208	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T19	vdd	I1/a2bar	I1/net1284	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T20	I1/net1284	I1/a1bar	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T14	I1/net160	I1/net1284	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T21	vdd	I1/a0bar	I1/net1284	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22U	PS=0.65U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI159/T2	vdd	I159/net32	I159/net28	vdd	pfet	L=0.12U
+ W=9.26U
+ AD=2.9632P	AS=2.9632P	PD=19.16U	PS=19.16U
+ wt=9.26e-06 wf=9.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.1352e-12 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0238741 nrd=0.0238741 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T591	vdd	addr0	I1/a0bar	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T592	vdd	addr1	I1/a1bar	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T23	I1/net156	addr0	vdd	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2376P	AS=0.2442P	PD=2.04U	PS=2.06U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.92e-14 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T50	I1/net144	addr1	vdd	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2376P	AS=0.2442P	PD=2.04U	PS=2.06U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.92e-14 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T22	I1/a0	I1/net156	vdd	vdd	pfet	L=0.12U	W=1.14U
+ AD=0.4104P	AS=0.4218P	PD=3U	PS=3.02U
+ wt=1.14e-06 wf=1.14e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=5.28e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.368e-13 nrs=0.200913 nrd=0.200913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T27	I1/a1	I1/net144	vdd	vdd	pfet	L=0.12U	W=1.14U
+ AD=0.4104P	AS=0.4218P	PD=3U	PS=3.02U
+ wt=1.14e-06 wf=1.14e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=5.82e-14 panw7=1.266e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=4.8e-15 nrs=0.200913 nrd=0.200913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI159/T0	vdd	clk	I159/net36	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=2.76e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.26e-14 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI159/T1	vdd	I159/net36	I159/net32	vdd	pfet	L=0.12U
+ W=2.48U
+ AD=0.7936P	AS=0.7936P	PD=5.6U	PS=5.6U
+ wt=2.48e-06 wf=2.48e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=3.216e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0903491 nrd=0.0903491 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T28	I1/a2	I1/net116	vdd	vdd	pfet	L=0.12U	W=1.14U
+ AD=0.4104P	AS=0.4218P	PD=3U	PS=3.02U
+ wt=1.14e-06 wf=1.14e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=5.82e-14 panw7=1.266e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=4.8e-15 nrs=0.200913 nrd=0.200913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3148/T1	I0/I3148/net13	I0/I3148/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3129/T1	I0/I3129/net13	I0/I3129/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3116/T0	vdd	I0/I3116/net13	I0/I3116/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3097/T0	vdd	I0/I3097/net13	I0/I3097/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3116/T1	I0/I3116/net13	I0/I3116/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3097/T1	I0/I3097/net13	I0/I3097/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3180/T0	vdd	I0/I3180/net13	I0/I3180/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3161/T0	vdd	I0/I3161/net13	I0/I3161/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3180/T1	I0/I3180/net13	I0/I3180/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3161/T1	I0/I3161/net13	I0/I3161/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3148/T0	vdd	I0/I3148/net13	I0/I3148/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3129/T0	vdd	I0/I3129/net13	I0/I3129/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I91/T1	I0/I91/net13	I0/I91/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I110/T1	I0/I110/net13	I0/I110/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3212/T0	vdd	I0/I3212/net13	I0/I3212/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3193/T0	vdd	I0/I3193/net13	I0/I3193/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3212/T1	I0/I3212/net13	I0/I3212/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3193/T1	I0/I3193/net13	I0/I3193/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3020/T0	vdd	I0/I3020/net13	I0/I3020/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3001/T0	vdd	I0/I3001/net13	I0/I3001/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3020/T1	I0/I3020/net13	I0/I3020/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3001/T1	I0/I3001/net13	I0/I3001/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I91/T0	vdd	I0/I91/net13	I0/I91/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I110/T0	vdd	I0/I110/net13	I0/I110/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3084/T1	I0/I3084/net13	I0/I3084/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3065/T1	I0/I3065/net13	I0/I3065/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3052/T0	vdd	I0/I3052/net13	I0/I3052/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3033/T0	vdd	I0/I3033/net13	I0/I3033/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3052/T1	I0/I3052/net13	I0/I3052/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3033/T1	I0/I3033/net13	I0/I3033/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I5/T0	vdd	I0/I5/net13	I0/I5/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2821/T0	vdd	I0/I2821/net13	I0/I2821/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I5/T1	I0/I5/net13	I0/I5/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2821/T1	I0/I2821/net13	I0/I2821/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3084/T0	vdd	I0/I3084/net13	I0/I3084/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3065/T0	vdd	I0/I3065/net13	I0/I3065/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2923/T1	I0/I2923/net13	I0/I2923/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2903/T1	I0/I2903/net13	I0/I2903/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2893/T0	vdd	I0/I2893/net13	I0/I2893/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2871/T0	vdd	I0/I2871/net13	I0/I2871/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2893/T1	I0/I2893/net13	I0/I2893/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2871/T1	I0/I2871/net13	I0/I2871/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2951/T0	vdd	I0/I2951/net13	I0/I2951/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2940/T0	vdd	I0/I2940/net13	I0/I2940/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2951/T1	I0/I2951/net13	I0/I2951/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.4e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.96e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2940/T1	I0/I2940/net13	I0/I2940/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.4e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.96e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2923/T0	vdd	I0/I2923/net13	I0/I2923/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2903/T0	vdd	I0/I2903/net13	I0/I2903/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T121	net952	I1/net1176	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T146	net951	I1/net1324	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T120	vdd	I1/net72	I1/net1176	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T119	I1/net1176	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T148	vdd	I1/net412	I1/net1324	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T147	I1/net1324	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T155	vdd	I1/net284	I1/net1492	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T117	vdd	I1/net160	I1/net1188	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T116	I1/net1188	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T115	vdd	I1/a4	I1/net1188	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T152	vdd	I1/net316	I1/net1420	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T151	I1/net1420	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T150	vdd	I1/a4bar	I1/net1420	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T158	vdd	I1/net316	I1/net1328	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T118	I1/net72	I1/net1188	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T149	I1/net412	I1/net1420	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T47	vdd	I1/net264	I1/net260	vdd	pfet	L=0.12U
+ W=1.65U
+ AD=0.6105P	AS=0.594P	PD=4.04U	PS=4.02U
+ wt=1.65e-06 wf=1.65e-06 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.64e-14 panw8=4.8e-14 panw7=2.256e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.137072 nrd=0.137072 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T593	vdd	addr2	I1/a2bar	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T53	I1/net116	addr2	vdd	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2376P	AS=0.2442P	PD=2.04U	PS=2.06U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.92e-14 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T153	I1/net316	I1/net1460	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T51	I1/a3	I1/net260	vdd	vdd	pfet	L=0.12U	W=4.1U
+ AD=1.476P	AS=1.517P	PD=8.92U	PS=8.94U
+ wt=4.1e-06 wf=4.1e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=5.196e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.054254 nrd=0.054254 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3144/T1	I0/I3144/net13	I0/I3144/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3142/T1	I0/I3142/net13	I0/I3142/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3138/T1	I0/I3138/net13	I0/I3138/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3112/T0	vdd	I0/I3112/net13	I0/I3112/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3110/T0	vdd	I0/I3110/net13	I0/I3110/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3106/T0	vdd	I0/I3106/net13	I0/I3106/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3112/T1	I0/I3112/net13	I0/I3112/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3110/T1	I0/I3110/net13	I0/I3110/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3106/T1	I0/I3106/net13	I0/I3106/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3176/T0	vdd	I0/I3176/net13	I0/I3176/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3174/T0	vdd	I0/I3174/net13	I0/I3174/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3170/T0	vdd	I0/I3170/net13	I0/I3170/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3176/T1	I0/I3176/net13	I0/I3176/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3174/T1	I0/I3174/net13	I0/I3174/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3170/T1	I0/I3170/net13	I0/I3170/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3144/T0	vdd	I0/I3144/net13	I0/I3144/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3142/T0	vdd	I0/I3142/net13	I0/I3142/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3138/T0	vdd	I0/I3138/net13	I0/I3138/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I95/T1	I0/I95/net13	I0/I95/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I97/T1	I0/I97/net13	I0/I97/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I101/T1	I0/I101/net13	I0/I101/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3208/T0	vdd	I0/I3208/net13	I0/I3208/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3206/T0	vdd	I0/I3206/net13	I0/I3206/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3202/T0	vdd	I0/I3202/net13	I0/I3202/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3208/T1	I0/I3208/net13	I0/I3208/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3206/T1	I0/I3206/net13	I0/I3206/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3202/T1	I0/I3202/net13	I0/I3202/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3016/T0	vdd	I0/I3016/net13	I0/I3016/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3014/T0	vdd	I0/I3014/net13	I0/I3014/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3010/T0	vdd	I0/I3010/net13	I0/I3010/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3016/T1	I0/I3016/net13	I0/I3016/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3014/T1	I0/I3014/net13	I0/I3014/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3010/T1	I0/I3010/net13	I0/I3010/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I95/T0	vdd	I0/I95/net13	I0/I95/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I97/T0	vdd	I0/I97/net13	I0/I97/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I101/T0	vdd	I0/I101/net13	I0/I101/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3080/T1	I0/I3080/net13	I0/I3080/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3078/T1	I0/I3078/net13	I0/I3078/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3074/T1	I0/I3074/net13	I0/I3074/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3048/T0	vdd	I0/I3048/net13	I0/I3048/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3046/T0	vdd	I0/I3046/net13	I0/I3046/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3042/T0	vdd	I0/I3042/net13	I0/I3042/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3048/T1	I0/I3048/net13	I0/I3048/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3046/T1	I0/I3046/net13	I0/I3046/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3042/T1	I0/I3042/net13	I0/I3042/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2812/T0	vdd	I0/I2812/net13	I0/I2812/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2825/T0	vdd	I0/I2825/net13	I0/I2825/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2805/T0	vdd	I0/I2805/net13	I0/I2805/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2812/T1	I0/I2812/net13	I0/I2812/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2825/T1	I0/I2825/net13	I0/I2825/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2805/T1	I0/I2805/net13	I0/I2805/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3080/T0	vdd	I0/I3080/net13	I0/I3080/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3078/T0	vdd	I0/I3078/net13	I0/I3078/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3074/T0	vdd	I0/I3074/net13	I0/I3074/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2922/T1	I0/I2922/net13	I0/I2922/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2919/T1	I0/I2919/net13	I0/I2919/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2910/T1	I0/I2910/net13	I0/I2910/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2877/T0	vdd	I0/I2877/net13	I0/I2877/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2879/T0	vdd	I0/I2879/net13	I0/I2879/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2886/T0	vdd	I0/I2886/net13	I0/I2886/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2877/T1	I0/I2877/net13	I0/I2877/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2879/T1	I0/I2879/net13	I0/I2879/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2886/T1	I0/I2886/net13	I0/I2886/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2956/T0	vdd	I0/I2956/net13	I0/I2956/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2957/T0	vdd	I0/I2957/net13	I0/I2957/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2936/T0	vdd	I0/I2936/net13	I0/I2936/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2956/T1	I0/I2956/net13	I0/I2956/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.96e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.4e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2957/T1	I0/I2957/net13	I0/I2957/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.96e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.4e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2936/T1	I0/I2936/net13	I0/I2936/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2922/T0	vdd	I0/I2922/net13	I0/I2922/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2919/T0	vdd	I0/I2919/net13	I0/I2919/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2910/T0	vdd	I0/I2910/net13	I0/I2910/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T156	I1/net1492	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T162	vdd	I1/net420	I1/net1436	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T163	I1/net1436	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T173	vdd	I1/net352	I1/net1452	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T172	I1/net1452	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T154	net950	I1/net1492	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T161	net949	I1/net1436	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T174	net948	I1/net1452	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T159	I1/net1328	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T160	vdd	I1/a4	I1/net1328	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T165	vdd	I1/net316	I1/net1496	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T166	I1/net1496	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T167	vdd	I1/a4bar	I1/net1496	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T170	vdd	I1/net316	I1/net1488	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T169	I1/net1488	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T168	vdd	I1/a4	I1/net1488	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T157	I1/net284	I1/net1328	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T164	I1/net420	I1/net1496	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T171	I1/net352	I1/net1488	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T143	vdd	I1/a2	I1/net1460	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T144	I1/net1460	I1/a1bar	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T145	vdd	I1/a0bar	I1/net1460	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22U	PS=0.65U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T40	I1/net264	I1/net124	vdd	vdd	pfet	L=0.12U
+ W=1.05U
+ AD=0.378P	AS=0.3885P	PD=2.82U	PS=2.84U
+ wt=1.05e-06 wf=1.05e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.2e-14 panw8=2.4e-14 panw7=1.5e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.218905 nrd=0.218905 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T36	vdd	addr3	I1/net124	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3098/T0	vdd	I0/I3098/net13	I0/I3098/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3099/T0	vdd	I0/I3099/net13	I0/I3099/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3089/T0	vdd	I0/I3089/net13	I0/I3089/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3115/T0	vdd	I0/I3115/net13	I0/I3115/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3109/T0	vdd	I0/I3109/net13	I0/I3109/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3098/T1	I0/I3098/net13	I0/I3098/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3099/T1	I0/I3099/net13	I0/I3099/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3089/T1	I0/I3089/net13	I0/I3089/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3115/T1	I0/I3115/net13	I0/I3115/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3109/T1	I0/I3109/net13	I0/I3109/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3130/T1	I0/I3130/net13	I0/I3130/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3131/T1	I0/I3131/net13	I0/I3131/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3121/T1	I0/I3121/net13	I0/I3121/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3147/T1	I0/I3147/net13	I0/I3147/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3141/T1	I0/I3141/net13	I0/I3141/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3130/T0	vdd	I0/I3130/net13	I0/I3130/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3131/T0	vdd	I0/I3131/net13	I0/I3131/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3121/T0	vdd	I0/I3121/net13	I0/I3121/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3147/T0	vdd	I0/I3147/net13	I0/I3147/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3141/T0	vdd	I0/I3141/net13	I0/I3141/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3162/T0	vdd	I0/I3162/net13	I0/I3162/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3163/T0	vdd	I0/I3163/net13	I0/I3163/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3153/T0	vdd	I0/I3153/net13	I0/I3153/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3179/T0	vdd	I0/I3179/net13	I0/I3179/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3173/T0	vdd	I0/I3173/net13	I0/I3173/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3162/T1	I0/I3162/net13	I0/I3162/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3163/T1	I0/I3163/net13	I0/I3163/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3153/T1	I0/I3153/net13	I0/I3153/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3179/T1	I0/I3179/net13	I0/I3179/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3173/T1	I0/I3173/net13	I0/I3173/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3194/T0	vdd	I0/I3194/net13	I0/I3194/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3195/T0	vdd	I0/I3195/net13	I0/I3195/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3185/T0	vdd	I0/I3185/net13	I0/I3185/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3211/T0	vdd	I0/I3211/net13	I0/I3211/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3205/T0	vdd	I0/I3205/net13	I0/I3205/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3194/T1	I0/I3194/net13	I0/I3194/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3195/T1	I0/I3195/net13	I0/I3195/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3185/T1	I0/I3185/net13	I0/I3185/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3211/T1	I0/I3211/net13	I0/I3211/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3205/T1	I0/I3205/net13	I0/I3205/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I109/T1	I0/I109/net13	I0/I109/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I108/T1	I0/I108/net13	I0/I108/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I118/T1	I0/I118/net13	I0/I118/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I92/T1	I0/I92/net13	I0/I92/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I98/T1	I0/I98/net13	I0/I98/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I109/T0	vdd	I0/I109/net13	I0/I109/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I108/T0	vdd	I0/I108/net13	I0/I108/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I118/T0	vdd	I0/I118/net13	I0/I118/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I92/T0	vdd	I0/I92/net13	I0/I92/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I98/T0	vdd	I0/I98/net13	I0/I98/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3002/T0	vdd	I0/I3002/net13	I0/I3002/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3003/T0	vdd	I0/I3003/net13	I0/I3003/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2993/T0	vdd	I0/I2993/net13	I0/I2993/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3019/T0	vdd	I0/I3019/net13	I0/I3019/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3013/T0	vdd	I0/I3013/net13	I0/I3013/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3002/T1	I0/I3002/net13	I0/I3002/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3003/T1	I0/I3003/net13	I0/I3003/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2993/T1	I0/I2993/net13	I0/I2993/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3019/T1	I0/I3019/net13	I0/I3019/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3013/T1	I0/I3013/net13	I0/I3013/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3034/T0	vdd	I0/I3034/net13	I0/I3034/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3035/T0	vdd	I0/I3035/net13	I0/I3035/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3025/T0	vdd	I0/I3025/net13	I0/I3025/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3051/T0	vdd	I0/I3051/net13	I0/I3051/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3045/T0	vdd	I0/I3045/net13	I0/I3045/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3034/T1	I0/I3034/net13	I0/I3034/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3035/T1	I0/I3035/net13	I0/I3035/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3025/T1	I0/I3025/net13	I0/I3025/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3051/T1	I0/I3051/net13	I0/I3051/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3045/T1	I0/I3045/net13	I0/I3045/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3066/T1	I0/I3066/net13	I0/I3066/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3067/T1	I0/I3067/net13	I0/I3067/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3057/T1	I0/I3057/net13	I0/I3057/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3083/T1	I0/I3083/net13	I0/I3083/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3077/T1	I0/I3077/net13	I0/I3077/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3066/T0	vdd	I0/I3066/net13	I0/I3066/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3067/T0	vdd	I0/I3067/net13	I0/I3067/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3057/T0	vdd	I0/I3057/net13	I0/I3057/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3083/T0	vdd	I0/I3083/net13	I0/I3083/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3077/T0	vdd	I0/I3077/net13	I0/I3077/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2826/T0	vdd	I0/I2826/net13	I0/I2826/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2816/T0	vdd	I0/I2816/net13	I0/I2816/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2803/T0	vdd	I0/I2803/net13	I0/I2803/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2811/T0	vdd	I0/I2811/net13	I0/I2811/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2813/T0	vdd	I0/I2813/net13	I0/I2813/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2826/T1	I0/I2826/net13	I0/I2826/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2816/T1	I0/I2816/net13	I0/I2816/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2803/T1	I0/I2803/net13	I0/I2803/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2811/T1	I0/I2811/net13	I0/I2811/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2813/T1	I0/I2813/net13	I0/I2813/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2872/T0	vdd	I0/I2872/net13	I0/I2872/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2887/T0	vdd	I0/I2887/net13	I0/I2887/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2889/T0	vdd	I0/I2889/net13	I0/I2889/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2880/T0	vdd	I0/I2880/net13	I0/I2880/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2881/T0	vdd	I0/I2881/net13	I0/I2881/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2872/T1	I0/I2872/net13	I0/I2872/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2887/T1	I0/I2887/net13	I0/I2887/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2889/T1	I0/I2889/net13	I0/I2889/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2880/T1	I0/I2880/net13	I0/I2880/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2881/T1	I0/I2881/net13	I0/I2881/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2905/T1	I0/I2905/net13	I0/I2905/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2920/T1	I0/I2920/net13	I0/I2920/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2915/T1	I0/I2915/net13	I0/I2915/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2902/T1	I0/I2902/net13	I0/I2902/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2901/T1	I0/I2901/net13	I0/I2901/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2905/T0	vdd	I0/I2905/net13	I0/I2905/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2920/T0	vdd	I0/I2920/net13	I0/I2920/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2915/T0	vdd	I0/I2915/net13	I0/I2915/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2902/T0	vdd	I0/I2902/net13	I0/I2902/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2901/T0	vdd	I0/I2901/net13	I0/I2901/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2941/T0	vdd	I0/I2941/net13	I0/I2941/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2953/T0	vdd	I0/I2953/net13	I0/I2953/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2949/T0	vdd	I0/I2949/net13	I0/I2949/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2938/T0	vdd	I0/I2938/net13	I0/I2938/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2935/T0	vdd	I0/I2935/net13	I0/I2935/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2941/T1	I0/I2941/net13	I0/I2941/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2953/T1	I0/I2953/net13	I0/I2953/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2949/T1	I0/I2949/net13	I0/I2949/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2938/T1	I0/I2938/net13	I0/I2938/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2935/T1	I0/I2935/net13	I0/I2935/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T235	net947	I1/net1644	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T227	net946	I1/net1616	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T220	net945	I1/net1588	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T207	net944	I1/net1544	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T233	vdd	I1/net532	I1/net1644	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T234	I1/net1644	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T226	vdd	I1/net492	I1/net1616	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T225	I1/net1616	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T219	vdd	I1/net456	I1/net1588	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T218	I1/net1588	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T208	vdd	I1/net452	I1/net1544	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T209	I1/net1544	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T276	vdd	I1/net600	I1/net1672	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T232	I1/net532	I1/net1628	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T224	I1/net492	I1/net1604	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T217	I1/net456	I1/net1576	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T210	I1/net452	I1/net1556	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T229	vdd	I1/net516	I1/net1628	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T230	I1/net1628	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T231	vdd	I1/a4bar	I1/net1628	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T223	vdd	I1/net516	I1/net1604	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T222	I1/net1604	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T221	vdd	I1/a4	I1/net1604	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T216	vdd	I1/net516	I1/net1576	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T215	I1/net1576	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T214	vdd	I1/a4bar	I1/net1576	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T211	vdd	I1/net516	I1/net1556	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T212	I1/net1556	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T213	vdd	I1/a4	I1/net1556	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T280	vdd	I1/net776	I1/net1840	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T68	vdd	addr3	I1/net328	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T49	vdd	I1/net212	I1/net256	vdd	pfet	L=0.12U
+ W=1.65U
+ AD=0.6105P	AS=0.594P	PD=4.04U	PS=4.02U
+ wt=1.65e-06 wf=1.65e-06 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=8.64e-14 panw8=4.8e-14 panw7=2.256e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.137072 nrd=0.137072 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T58	I1/net320	I1/net328	vdd	vdd	pfet	L=0.12U
+ W=1.65U
+ AD=0.594P	AS=0.6105P	PD=4.02U	PS=4.04U
+ wt=1.65e-06 wf=1.65e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.22e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=6.6e-14 nrs=0.137072 nrd=0.137072 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T57	I1/a3bar	I1/net320	vdd	vdd	pfet	L=0.12U
+ W=4.1U
+ AD=1.476P	AS=1.517P	PD=8.92U	PS=8.94U
+ wt=4.1e-06 wf=4.1e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=5.196e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.054254 nrd=0.054254 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T238	vdd	I1/a2bar	I1/net1656	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T237	I1/net1656	I1/a1	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T228	I1/net516	I1/net1656	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T236	vdd	I1/a0bar	I1/net1656	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22U	PS=0.65U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T52	I1/a4	I1/net256	vdd	vdd	pfet	L=0.12U	W=4.1U
+ AD=1.476P	AS=1.517P	PD=8.92U	PS=8.94U
+ wt=4.1e-06 wf=4.1e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=5.196e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.054254 nrd=0.054254 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3127/T1	I0/I3127/net13	I0/I3127/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3120/T1	I0/I3120/net13	I0/I3120/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3095/T0	vdd	I0/I3095/net13	I0/I3095/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3088/T0	vdd	I0/I3088/net13	I0/I3088/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3095/T1	I0/I3095/net13	I0/I3095/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3088/T1	I0/I3088/net13	I0/I3088/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3159/T0	vdd	I0/I3159/net13	I0/I3159/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3152/T0	vdd	I0/I3152/net13	I0/I3152/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3159/T1	I0/I3159/net13	I0/I3159/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3152/T1	I0/I3152/net13	I0/I3152/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3127/T0	vdd	I0/I3127/net13	I0/I3127/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3120/T0	vdd	I0/I3120/net13	I0/I3120/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I112/T1	I0/I112/net13	I0/I112/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I119/T1	I0/I119/net13	I0/I119/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3191/T0	vdd	I0/I3191/net13	I0/I3191/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3184/T0	vdd	I0/I3184/net13	I0/I3184/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3191/T1	I0/I3191/net13	I0/I3191/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3184/T1	I0/I3184/net13	I0/I3184/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2999/T0	vdd	I0/I2999/net13	I0/I2999/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2992/T0	vdd	I0/I2992/net13	I0/I2992/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2999/T1	I0/I2999/net13	I0/I2999/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2992/T1	I0/I2992/net13	I0/I2992/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I112/T0	vdd	I0/I112/net13	I0/I112/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I119/T0	vdd	I0/I119/net13	I0/I119/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3063/T1	I0/I3063/net13	I0/I3063/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3056/T1	I0/I3056/net13	I0/I3056/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3031/T0	vdd	I0/I3031/net13	I0/I3031/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3024/T0	vdd	I0/I3024/net13	I0/I3024/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3031/T1	I0/I3031/net13	I0/I3031/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3024/T1	I0/I3024/net13	I0/I3024/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2827/T0	vdd	I0/I2827/net13	I0/I2827/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2804/T0	vdd	I0/I2804/net13	I0/I2804/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2827/T1	I0/I2827/net13	I0/I2827/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2804/T1	I0/I2804/net13	I0/I2804/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3063/T0	vdd	I0/I3063/net13	I0/I3063/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3056/T0	vdd	I0/I3056/net13	I0/I3056/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2914/T1	I0/I2914/net13	I0/I2914/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2913/T1	I0/I2913/net13	I0/I2913/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2865/T0	vdd	I0/I2865/net13	I0/I2865/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2890/T0	vdd	I0/I2890/net13	I0/I2890/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2865/T1	I0/I2865/net13	I0/I2865/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2890/T1	I0/I2890/net13	I0/I2890/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2947/T0	vdd	I0/I2947/net13	I0/I2947/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2950/T0	vdd	I0/I2950/net13	I0/I2950/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2947/T1	I0/I2947/net13	I0/I2947/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2950/T1	I0/I2950/net13	I0/I2950/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2914/T0	vdd	I0/I2914/net13	I0/I2914/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2913/T0	vdd	I0/I2913/net13	I0/I2913/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T275	I1/net1672	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T283	vdd	I1/net768	I1/net1464	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T284	I1/net1464	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T290	vdd	I1/net704	I1/net1816	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T291	I1/net1816	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T274	net943	I1/net1672	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T282	net942	I1/net1464	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T289	net941	I1/net1816	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T279	I1/net1840	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T278	vdd	I1/a4bar	I1/net1840	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T286	vdd	I1/net776	I1/net1792	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T287	I1/net1792	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T288	vdd	I1/a4	I1/net1792	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T293	vdd	I1/net776	I1/net1352	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T294	I1/net1352	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T277	I1/net600	I1/net1840	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T285	I1/net768	I1/net1792	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T292	I1/net704	I1/net1352	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T271	vdd	I1/a2	I1/net1820	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T272	I1/net1820	I1/a1	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T281	I1/net776	I1/net1820	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T273	vdd	I1/a0bar	I1/net1820	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22U	PS=0.65U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T42	I1/net212	I1/net120	vdd	vdd	pfet	L=0.12U
+ W=1.05U
+ AD=0.378P	AS=0.3885P	PD=2.82U	PS=2.84U
+ wt=1.05e-06 wf=1.05e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.2e-14 panw8=2.4e-14 panw7=1.5e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.218905 nrd=0.218905 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T39	vdd	addr4	I1/net120	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T295	vdd	I1/a4bar	I1/net1352	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3175/T0	vdd	I0/I3175/net13	I0/I3175/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3175/T1	I0/I3175/net13	I0/I3175/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3143/T0	vdd	I0/I3143/net13	I0/I3143/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3143/T1	I0/I3143/net13	I0/I3143/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3111/T0	vdd	I0/I3111/net13	I0/I3111/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3111/T1	I0/I3111/net13	I0/I3111/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3015/T0	vdd	I0/I3015/net13	I0/I3015/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3015/T1	I0/I3015/net13	I0/I3015/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I96/T0	vdd	I0/I96/net13	I0/I96/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I96/T1	I0/I96/net13	I0/I96/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3207/T0	vdd	I0/I3207/net13	I0/I3207/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3207/T1	I0/I3207/net13	I0/I3207/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2802/T0	vdd	I0/I2802/net13	I0/I2802/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2802/T1	I0/I2802/net13	I0/I2802/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3079/T0	vdd	I0/I3079/net13	I0/I3079/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3079/T1	I0/I3079/net13	I0/I3079/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3047/T0	vdd	I0/I3047/net13	I0/I3047/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3047/T1	I0/I3047/net13	I0/I3047/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2943/T0	vdd	I0/I2943/net13	I0/I2943/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2943/T1	I0/I2943/net13	I0/I2943/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2908/T0	vdd	I0/I2908/net13	I0/I2908/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2908/T1	I0/I2908/net13	I0/I2908/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2891/T0	vdd	I0/I2891/net13	I0/I2891/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2891/T1	I0/I2891/net13	I0/I2891/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T298	vdd	I1/net776	I1/net1880	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T297	I1/net1880	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T299	I1/net708	I1/net1880	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T301	vdd	I1/net708	I1/net1852	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T300	I1/net1852	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T302	net940	I1/net1852	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T296	vdd	I1/a4	I1/net1880	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI0/I3172/T0	vdd	I0/I3172/net13	I0/I3172/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3172/T1	I0/I3172/net13	I0/I3172/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3140/T0	vdd	I0/I3140/net13	I0/I3140/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3140/T1	I0/I3140/net13	I0/I3140/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3108/T0	vdd	I0/I3108/net13	I0/I3108/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3108/T1	I0/I3108/net13	I0/I3108/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3012/T0	vdd	I0/I3012/net13	I0/I3012/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3012/T1	I0/I3012/net13	I0/I3012/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I99/T0	vdd	I0/I99/net13	I0/I99/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I99/T1	I0/I99/net13	I0/I99/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3204/T0	vdd	I0/I3204/net13	I0/I3204/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3204/T1	I0/I3204/net13	I0/I3204/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2820/T0	vdd	I0/I2820/net13	I0/I2820/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2820/T1	I0/I2820/net13	I0/I2820/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3076/T0	vdd	I0/I3076/net13	I0/I3076/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3076/T1	I0/I3076/net13	I0/I3076/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3044/T0	vdd	I0/I3044/net13	I0/I3044/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3044/T1	I0/I3044/net13	I0/I3044/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2948/T0	vdd	I0/I2948/net13	I0/I2948/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2948/T1	I0/I2948/net13	I0/I2948/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2912/T0	vdd	I0/I2912/net13	I0/I2912/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2912/T1	I0/I2912/net13	I0/I2912/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2875/T0	vdd	I0/I2875/net13	I0/I2875/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2875/T1	I0/I2875/net13	I0/I2875/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T363	net939	I1/net1904	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T86	vdd	addr4	I1/net216	vdd	pfet	L=0.12U	W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.92e-14 panw7=1.032e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T357	vdd	I1/net616	I1/net1716	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T358	I1/net1716	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T359	vdd	I1/a4bar	I1/net1716	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T360	I1/net788	I1/net1716	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96U	PS=2.98U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T361	vdd	I1/net788	I1/net1904	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T362	I1/net1904	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T70	I1/net336	I1/net216	vdd	vdd	pfet	L=0.12U
+ W=1.65U
+ AD=0.594P	AS=0.6105P	PD=4.02U	PS=4.04U
+ wt=1.65e-06 wf=1.65e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.22e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=6.6e-14 nrs=0.137072 nrd=0.137072 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T85	I1/a4bar	I1/net336	vdd	vdd	pfet	L=0.12U
+ W=4.1U
+ AD=1.476P	AS=1.517P	PD=8.92U	PS=8.94U
+ wt=4.1e-06 wf=4.1e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=5.196e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.054254 nrd=0.054254 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T356	I1/net616	I1/net1860	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3086/T1	I0/I3086/net13	I0/I3086/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3087/T1	I0/I3087/net13	I0/I3087/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3094/T1	I0/I3094/net13	I0/I3094/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3096/T1	I0/I3096/net13	I0/I3096/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3102/T1	I0/I3102/net13	I0/I3102/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3104/T1	I0/I3104/net13	I0/I3104/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3093/T1	I0/I3093/net13	I0/I3093/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3107/T1	I0/I3107/net13	I0/I3107/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3101/T1	I0/I3101/net13	I0/I3101/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3105/T1	I0/I3105/net13	I0/I3105/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3086/T0	vdd	I0/I3086/net13	I0/I3086/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3087/T0	vdd	I0/I3087/net13	I0/I3087/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3094/T0	vdd	I0/I3094/net13	I0/I3094/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3096/T0	vdd	I0/I3096/net13	I0/I3096/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3102/T0	vdd	I0/I3102/net13	I0/I3102/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3104/T0	vdd	I0/I3104/net13	I0/I3104/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3093/T0	vdd	I0/I3093/net13	I0/I3093/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3107/T0	vdd	I0/I3107/net13	I0/I3107/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3101/T0	vdd	I0/I3101/net13	I0/I3101/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3105/T0	vdd	I0/I3105/net13	I0/I3105/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3118/T1	I0/I3118/net13	I0/I3118/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3119/T1	I0/I3119/net13	I0/I3119/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3126/T1	I0/I3126/net13	I0/I3126/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3128/T1	I0/I3128/net13	I0/I3128/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3134/T1	I0/I3134/net13	I0/I3134/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3136/T1	I0/I3136/net13	I0/I3136/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3125/T1	I0/I3125/net13	I0/I3125/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3139/T1	I0/I3139/net13	I0/I3139/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3133/T1	I0/I3133/net13	I0/I3133/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3137/T1	I0/I3137/net13	I0/I3137/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3118/T0	vdd	I0/I3118/net13	I0/I3118/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3119/T0	vdd	I0/I3119/net13	I0/I3119/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3126/T0	vdd	I0/I3126/net13	I0/I3126/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3128/T0	vdd	I0/I3128/net13	I0/I3128/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3134/T0	vdd	I0/I3134/net13	I0/I3134/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3136/T0	vdd	I0/I3136/net13	I0/I3136/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3125/T0	vdd	I0/I3125/net13	I0/I3125/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3139/T0	vdd	I0/I3139/net13	I0/I3139/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3133/T0	vdd	I0/I3133/net13	I0/I3133/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3137/T0	vdd	I0/I3137/net13	I0/I3137/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3150/T1	I0/I3150/net13	I0/I3150/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3151/T1	I0/I3151/net13	I0/I3151/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3158/T1	I0/I3158/net13	I0/I3158/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3160/T1	I0/I3160/net13	I0/I3160/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3166/T1	I0/I3166/net13	I0/I3166/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3168/T1	I0/I3168/net13	I0/I3168/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3157/T1	I0/I3157/net13	I0/I3157/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3171/T1	I0/I3171/net13	I0/I3171/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3165/T1	I0/I3165/net13	I0/I3165/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3169/T1	I0/I3169/net13	I0/I3169/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3150/T0	vdd	I0/I3150/net13	I0/I3150/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3151/T0	vdd	I0/I3151/net13	I0/I3151/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3158/T0	vdd	I0/I3158/net13	I0/I3158/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3160/T0	vdd	I0/I3160/net13	I0/I3160/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3166/T0	vdd	I0/I3166/net13	I0/I3166/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3168/T0	vdd	I0/I3168/net13	I0/I3168/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3157/T0	vdd	I0/I3157/net13	I0/I3157/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3171/T0	vdd	I0/I3171/net13	I0/I3171/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3165/T0	vdd	I0/I3165/net13	I0/I3165/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3169/T0	vdd	I0/I3169/net13	I0/I3169/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3182/T1	I0/I3182/net13	I0/I3182/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3183/T1	I0/I3183/net13	I0/I3183/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3190/T1	I0/I3190/net13	I0/I3190/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3192/T1	I0/I3192/net13	I0/I3192/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3198/T1	I0/I3198/net13	I0/I3198/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3200/T1	I0/I3200/net13	I0/I3200/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3189/T1	I0/I3189/net13	I0/I3189/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3203/T1	I0/I3203/net13	I0/I3203/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3197/T1	I0/I3197/net13	I0/I3197/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3201/T1	I0/I3201/net13	I0/I3201/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3182/T0	vdd	I0/I3182/net13	I0/I3182/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3183/T0	vdd	I0/I3183/net13	I0/I3183/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3190/T0	vdd	I0/I3190/net13	I0/I3190/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3192/T0	vdd	I0/I3192/net13	I0/I3192/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3198/T0	vdd	I0/I3198/net13	I0/I3198/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3200/T0	vdd	I0/I3200/net13	I0/I3200/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3189/T0	vdd	I0/I3189/net13	I0/I3189/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3203/T0	vdd	I0/I3203/net13	I0/I3203/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3197/T0	vdd	I0/I3197/net13	I0/I3197/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3201/T0	vdd	I0/I3201/net13	I0/I3201/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I121/T1	I0/I121/net13	I0/I121/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I120/T1	I0/I120/net13	I0/I120/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I113/T1	I0/I113/net13	I0/I113/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I111/T1	I0/I111/net13	I0/I111/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I105/T1	I0/I105/net13	I0/I105/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I103/T1	I0/I103/net13	I0/I103/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I114/T1	I0/I114/net13	I0/I114/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I100/T1	I0/I100/net13	I0/I100/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I106/T1	I0/I106/net13	I0/I106/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I102/T1	I0/I102/net13	I0/I102/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I121/T0	vdd	I0/I121/net13	I0/I121/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I120/T0	vdd	I0/I120/net13	I0/I120/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I113/T0	vdd	I0/I113/net13	I0/I113/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I111/T0	vdd	I0/I111/net13	I0/I111/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I105/T0	vdd	I0/I105/net13	I0/I105/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I103/T0	vdd	I0/I103/net13	I0/I103/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I114/T0	vdd	I0/I114/net13	I0/I114/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I100/T0	vdd	I0/I100/net13	I0/I100/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I106/T0	vdd	I0/I106/net13	I0/I106/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I102/T0	vdd	I0/I102/net13	I0/I102/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2990/T1	I0/I2990/net13	I0/I2990/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2991/T1	I0/I2991/net13	I0/I2991/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2998/T1	I0/I2998/net13	I0/I2998/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3000/T1	I0/I3000/net13	I0/I3000/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3006/T1	I0/I3006/net13	I0/I3006/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3008/T1	I0/I3008/net13	I0/I3008/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2997/T1	I0/I2997/net13	I0/I2997/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3011/T1	I0/I3011/net13	I0/I3011/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3005/T1	I0/I3005/net13	I0/I3005/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3009/T1	I0/I3009/net13	I0/I3009/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2990/T0	vdd	I0/I2990/net13	I0/I2990/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2991/T0	vdd	I0/I2991/net13	I0/I2991/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2998/T0	vdd	I0/I2998/net13	I0/I2998/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3000/T0	vdd	I0/I3000/net13	I0/I3000/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3006/T0	vdd	I0/I3006/net13	I0/I3006/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3008/T0	vdd	I0/I3008/net13	I0/I3008/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2997/T0	vdd	I0/I2997/net13	I0/I2997/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3011/T0	vdd	I0/I3011/net13	I0/I3011/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3005/T0	vdd	I0/I3005/net13	I0/I3005/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3009/T0	vdd	I0/I3009/net13	I0/I3009/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3022/T1	I0/I3022/net13	I0/I3022/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3023/T1	I0/I3023/net13	I0/I3023/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3030/T1	I0/I3030/net13	I0/I3030/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3032/T1	I0/I3032/net13	I0/I3032/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3038/T1	I0/I3038/net13	I0/I3038/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3040/T1	I0/I3040/net13	I0/I3040/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3029/T1	I0/I3029/net13	I0/I3029/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3043/T1	I0/I3043/net13	I0/I3043/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3037/T1	I0/I3037/net13	I0/I3037/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3041/T1	I0/I3041/net13	I0/I3041/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3022/T0	vdd	I0/I3022/net13	I0/I3022/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3023/T0	vdd	I0/I3023/net13	I0/I3023/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3030/T0	vdd	I0/I3030/net13	I0/I3030/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3032/T0	vdd	I0/I3032/net13	I0/I3032/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3038/T0	vdd	I0/I3038/net13	I0/I3038/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3040/T0	vdd	I0/I3040/net13	I0/I3040/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3029/T0	vdd	I0/I3029/net13	I0/I3029/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3043/T0	vdd	I0/I3043/net13	I0/I3043/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3037/T0	vdd	I0/I3037/net13	I0/I3037/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3041/T0	vdd	I0/I3041/net13	I0/I3041/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3054/T1	I0/I3054/net13	I0/I3054/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3055/T1	I0/I3055/net13	I0/I3055/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3062/T1	I0/I3062/net13	I0/I3062/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3064/T1	I0/I3064/net13	I0/I3064/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3070/T1	I0/I3070/net13	I0/I3070/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3072/T1	I0/I3072/net13	I0/I3072/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3061/T1	I0/I3061/net13	I0/I3061/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3075/T1	I0/I3075/net13	I0/I3075/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3069/T1	I0/I3069/net13	I0/I3069/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3073/T1	I0/I3073/net13	I0/I3073/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3054/T0	vdd	I0/I3054/net13	I0/I3054/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3055/T0	vdd	I0/I3055/net13	I0/I3055/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3062/T0	vdd	I0/I3062/net13	I0/I3062/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3064/T0	vdd	I0/I3064/net13	I0/I3064/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3070/T0	vdd	I0/I3070/net13	I0/I3070/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3072/T0	vdd	I0/I3072/net13	I0/I3072/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3061/T0	vdd	I0/I3061/net13	I0/I3061/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3075/T0	vdd	I0/I3075/net13	I0/I3075/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3069/T0	vdd	I0/I3069/net13	I0/I3069/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3073/T0	vdd	I0/I3073/net13	I0/I3073/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2800/T1	I0/I2800/net13	I0/I2800/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2810/T1	I0/I2810/net13	I0/I2810/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2809/T1	I0/I2809/net13	I0/I2809/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2801/T1	I0/I2801/net13	I0/I2801/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2823/T1	I0/I2823/net13	I0/I2823/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2824/T1	I0/I2824/net13	I0/I2824/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2808/T1	I0/I2808/net13	I0/I2808/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2819/T1	I0/I2819/net13	I0/I2819/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2815/T1	I0/I2815/net13	I0/I2815/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2814/T1	I0/I2814/net13	I0/I2814/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2800/T0	vdd	I0/I2800/net13	I0/I2800/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2810/T0	vdd	I0/I2810/net13	I0/I2810/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2809/T0	vdd	I0/I2809/net13	I0/I2809/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2801/T0	vdd	I0/I2801/net13	I0/I2801/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2823/T0	vdd	I0/I2823/net13	I0/I2823/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2824/T0	vdd	I0/I2824/net13	I0/I2824/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2808/T0	vdd	I0/I2808/net13	I0/I2808/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2819/T0	vdd	I0/I2819/net13	I0/I2819/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2815/T0	vdd	I0/I2815/net13	I0/I2815/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2814/T0	vdd	I0/I2814/net13	I0/I2814/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2883/T1	I0/I2883/net13	I0/I2883/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2885/T1	I0/I2885/net13	I0/I2885/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2864/T1	I0/I2864/net13	I0/I2864/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2867/T1	I0/I2867/net13	I0/I2867/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2868/T1	I0/I2868/net13	I0/I2868/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2874/T1	I0/I2874/net13	I0/I2874/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2892/T1	I0/I2892/net13	I0/I2892/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2882/T1	I0/I2882/net13	I0/I2882/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2873/T1	I0/I2873/net13	I0/I2873/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2876/T1	I0/I2876/net13	I0/I2876/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2883/T0	vdd	I0/I2883/net13	I0/I2883/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2885/T0	vdd	I0/I2885/net13	I0/I2885/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2864/T0	vdd	I0/I2864/net13	I0/I2864/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2867/T0	vdd	I0/I2867/net13	I0/I2867/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2868/T0	vdd	I0/I2868/net13	I0/I2868/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2874/T0	vdd	I0/I2874/net13	I0/I2874/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2892/T0	vdd	I0/I2892/net13	I0/I2892/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2882/T0	vdd	I0/I2882/net13	I0/I2882/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2873/T0	vdd	I0/I2873/net13	I0/I2873/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2876/T0	vdd	I0/I2876/net13	I0/I2876/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2918/T1	I0/I2918/net13	I0/I2918/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2906/T1	I0/I2906/net13	I0/I2906/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2916/T1	I0/I2916/net13	I0/I2916/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2896/T1	I0/I2896/net13	I0/I2896/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2897/T1	I0/I2897/net13	I0/I2897/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2907/T1	I0/I2907/net13	I0/I2907/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2917/T1	I0/I2917/net13	I0/I2917/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2924/T1	I0/I2924/net13	I0/I2924/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2921/T1	I0/I2921/net13	I0/I2921/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2911/T1	I0/I2911/net13	I0/I2911/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2918/T0	vdd	I0/I2918/net13	I0/I2918/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2906/T0	vdd	I0/I2906/net13	I0/I2906/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2916/T0	vdd	I0/I2916/net13	I0/I2916/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2896/T0	vdd	I0/I2896/net13	I0/I2896/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2897/T0	vdd	I0/I2897/net13	I0/I2897/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2907/T0	vdd	I0/I2907/net13	I0/I2907/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2917/T0	vdd	I0/I2917/net13	I0/I2917/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2924/T0	vdd	I0/I2924/net13	I0/I2924/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2921/T0	vdd	I0/I2921/net13	I0/I2921/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2911/T0	vdd	I0/I2911/net13	I0/I2911/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2952/T1	I0/I2952/net13	I0/I2952/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2942/T1	I0/I2942/net13	I0/I2942/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2932/T1	I0/I2932/net13	I0/I2932/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2928/T1	I0/I2928/net13	I0/I2928/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2929/T1	I0/I2929/net13	I0/I2929/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2945/T1	I0/I2945/net13	I0/I2945/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2954/T1	I0/I2954/net13	I0/I2954/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2955/T1	I0/I2955/net13	I0/I2955/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2946/T1	I0/I2946/net13	I0/I2946/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2944/T1	I0/I2944/net13	I0/I2944/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2952/T0	vdd	I0/I2952/net13	I0/I2952/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2942/T0	vdd	I0/I2942/net13	I0/I2942/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2932/T0	vdd	I0/I2932/net13	I0/I2932/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2928/T0	vdd	I0/I2928/net13	I0/I2928/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2929/T0	vdd	I0/I2929/net13	I0/I2929/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2945/T0	vdd	I0/I2945/net13	I0/I2945/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2954/T0	vdd	I0/I2954/net13	I0/I2954/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2955/T0	vdd	I0/I2955/net13	I0/I2955/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2946/T0	vdd	I0/I2946/net13	I0/I2946/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2944/T0	vdd	I0/I2944/net13	I0/I2944/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T354	vdd	I1/net796	I1/net1772	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T353	I1/net1772	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T347	vdd	I1/net732	I1/net1752	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T346	I1/net1752	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T336	vdd	I1/net812	I1/net1708	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T355	net938	I1/net1772	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T348	net937	I1/net1752	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T337	I1/net1708	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T404	vdd	I1/net864	I1/net1944	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T403	I1/net1944	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T411	vdd	I1/net908	I1/net1972	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T335	net936	I1/net1708	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T402	net935	I1/net1944	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T412	I1/net1972	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T418	vdd	I1/net944	I1/net2000	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T419	I1/net2000	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T429	vdd	I1/net948	I1/net2044	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T428	I1/net2044	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T410	net934	I1/net1972	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T417	net933	I1/net2000	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T430	net932	I1/net2044	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T489	vdd	I1/net1076	I1/net2096	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T490	I1/net2096	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T482	vdd	I1/net1116	I1/net2140	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T481	I1/net2140	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T491	net931	I1/net2096	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T483	net930	I1/net2140	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T352	I1/net796	I1/net1800	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T345	I1/net732	I1/net1780	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T338	I1/net812	I1/net1484	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T405	I1/net864	I1/net1960	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T413	I1/net908	I1/net1984	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T420	I1/net944	I1/net2012	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T427	I1/net948	I1/net2032	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T488	I1/net1076	I1/net1908	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T480	I1/net1116	I1/net1396	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T351	vdd	I1/net616	I1/net1800	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T350	I1/net1800	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T349	vdd	I1/a4	I1/net1800	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T344	vdd	I1/net616	I1/net1780	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T343	I1/net1780	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T342	vdd	I1/a4bar	I1/net1780	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T339	vdd	I1/net616	I1/net1484	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T340	I1/net1484	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T341	vdd	I1/a4	I1/net1484	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T408	vdd	I1/net880	I1/net1960	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T407	I1/net1960	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T406	vdd	I1/a4bar	I1/net1960	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T414	vdd	I1/net880	I1/net1984	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T415	I1/net1984	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T416	vdd	I1/a4	I1/net1984	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T421	vdd	I1/net880	I1/net2012	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T422	I1/net2012	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T423	vdd	I1/a4bar	I1/net2012	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T426	vdd	I1/net880	I1/net2032	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T425	I1/net2032	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T424	vdd	I1/a4	I1/net2032	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T485	vdd	I1/net1056	I1/net1908	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T486	I1/net1908	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T487	vdd	I1/a4bar	I1/net1908	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T479	vdd	I1/net1056	I1/net1396	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.4U	PS=0.74U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T478	I1/net1396	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74U	PS=0.75U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T477	vdd	I1/a4	I1/net1396	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75U	PS=1.4U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T364	vdd	I1/a0	I1/net1860	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22001U	PS=0.65001U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T401	vdd	I1/a0	I1/net1932	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22001U	PS=0.65001U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T492	vdd	I1/a0	I1/net2136	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22001U	PS=0.65001U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T38	vdd	addr_en	I1/net02041	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2442P	AS=0.2376P	PD=2.06U	PS=2.04U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=1.56e-14 panw7=1.068e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T35	vdd	I1/net02030	I1/net02033	vdd	pfet	L=0.12U
+ W=8.39U
+ AD=3.1043P	AS=3.0204P	PD=17.52U	PS=17.5U
+ wt=8.39e-06 wf=8.39e-06 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.0308e-12 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0263631 nrd=0.0263631 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T37	I1/net02030	I1/net02041	vdd	vdd	pfet	L=0.12U
+ W=2.36U
+ AD=0.8496P	AS=0.8732P	PD=5.44U	PS=5.46U
+ wt=2.36e-06 wf=2.36e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=3.072e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0950324 nrd=0.0950324 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T366	vdd	I1/a2bar	I1/net1860	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T399	vdd	I1/a2	I1/net1932	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T494	vdd	I1/a2bar	I1/net2136	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66U	PS=1.22U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T365	I1/net1860	I1/a1bar	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T400	I1/net1932	I1/a1bar	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T493	I1/net2136	I1/a1	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65U	PS=0.66U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T409	I1/net880	I1/net1932	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T484	I1/net1056	I1/net2136	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44U	PS=2.46U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T30	vdd	I1/net02033	I1/addr_en_b	vdd	pfet	L=0.12U
+ W=29.7U
+ AD=10.989P	AS=10.692P	PD=60.14U	PS=60.12U
+ wt=2.97e-05 wf=2.97e-05 sd=0 sb=3.7e-07 sa=3.6e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=3.5916e-12 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.00741865 nrd=0.00741865 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3117/T0	vdd	I0/I3117/net13	I0/I3117/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3103/T0	vdd	I0/I3103/net13	I0/I3103/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3114/T0	vdd	I0/I3114/net13	I0/I3114/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3113/T0	vdd	I0/I3113/net13	I0/I3113/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3090/T0	vdd	I0/I3090/net13	I0/I3090/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3117/T1	I0/I3117/net13	I0/I3117/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3103/T1	I0/I3103/net13	I0/I3103/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3114/T1	I0/I3114/net13	I0/I3114/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3113/T1	I0/I3113/net13	I0/I3113/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3090/T1	I0/I3090/net13	I0/I3090/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3149/T1	I0/I3149/net13	I0/I3149/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3135/T1	I0/I3135/net13	I0/I3135/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3146/T1	I0/I3146/net13	I0/I3146/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3145/T1	I0/I3145/net13	I0/I3145/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3122/T1	I0/I3122/net13	I0/I3122/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3149/T0	vdd	I0/I3149/net13	I0/I3149/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3135/T0	vdd	I0/I3135/net13	I0/I3135/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3146/T0	vdd	I0/I3146/net13	I0/I3146/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3145/T0	vdd	I0/I3145/net13	I0/I3145/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3122/T0	vdd	I0/I3122/net13	I0/I3122/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3181/T0	vdd	I0/I3181/net13	I0/I3181/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3167/T0	vdd	I0/I3167/net13	I0/I3167/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3178/T0	vdd	I0/I3178/net13	I0/I3178/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3177/T0	vdd	I0/I3177/net13	I0/I3177/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3154/T0	vdd	I0/I3154/net13	I0/I3154/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3181/T1	I0/I3181/net13	I0/I3181/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3167/T1	I0/I3167/net13	I0/I3167/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3178/T1	I0/I3178/net13	I0/I3178/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3177/T1	I0/I3177/net13	I0/I3177/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3154/T1	I0/I3154/net13	I0/I3154/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3213/T0	vdd	I0/I3213/net13	I0/I3213/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3199/T0	vdd	I0/I3199/net13	I0/I3199/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3210/T0	vdd	I0/I3210/net13	I0/I3210/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3209/T0	vdd	I0/I3209/net13	I0/I3209/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3186/T0	vdd	I0/I3186/net13	I0/I3186/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3213/T1	I0/I3213/net13	I0/I3213/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3199/T1	I0/I3199/net13	I0/I3199/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3210/T1	I0/I3210/net13	I0/I3210/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3209/T1	I0/I3209/net13	I0/I3209/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3186/T1	I0/I3186/net13	I0/I3186/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I90/T1	I0/I90/net13	I0/I90/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I104/T1	I0/I104/net13	I0/I104/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I93/T1	I0/I93/net13	I0/I93/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I94/T1	I0/I94/net13	I0/I94/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I117/T1	I0/I117/net13	I0/I117/net049	vdd	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I90/T0	vdd	I0/I90/net13	I0/I90/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I104/T0	vdd	I0/I104/net13	I0/I104/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I93/T0	vdd	I0/I93/net13	I0/I93/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I94/T0	vdd	I0/I94/net13	I0/I94/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I117/T0	vdd	I0/I117/net13	I0/I117/net049	vdd	pfet	L=0.12U
+ W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3021/T0	vdd	I0/I3021/net13	I0/I3021/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3007/T0	vdd	I0/I3007/net13	I0/I3007/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3018/T0	vdd	I0/I3018/net13	I0/I3018/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3017/T0	vdd	I0/I3017/net13	I0/I3017/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2994/T0	vdd	I0/I2994/net13	I0/I2994/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3021/T1	I0/I3021/net13	I0/I3021/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3007/T1	I0/I3007/net13	I0/I3007/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3018/T1	I0/I3018/net13	I0/I3018/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3017/T1	I0/I3017/net13	I0/I3017/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2994/T1	I0/I2994/net13	I0/I2994/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3053/T0	vdd	I0/I3053/net13	I0/I3053/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3039/T0	vdd	I0/I3039/net13	I0/I3039/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3050/T0	vdd	I0/I3050/net13	I0/I3050/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3049/T0	vdd	I0/I3049/net13	I0/I3049/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3026/T0	vdd	I0/I3026/net13	I0/I3026/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3053/T1	I0/I3053/net13	I0/I3053/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3039/T1	I0/I3039/net13	I0/I3039/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3050/T1	I0/I3050/net13	I0/I3050/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3049/T1	I0/I3049/net13	I0/I3049/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3026/T1	I0/I3026/net13	I0/I3026/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3085/T1	I0/I3085/net13	I0/I3085/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3071/T1	I0/I3071/net13	I0/I3071/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3082/T1	I0/I3082/net13	I0/I3082/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3081/T1	I0/I3081/net13	I0/I3081/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3058/T1	I0/I3058/net13	I0/I3058/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3085/T0	vdd	I0/I3085/net13	I0/I3085/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3071/T0	vdd	I0/I3071/net13	I0/I3071/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3082/T0	vdd	I0/I3082/net13	I0/I3082/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3081/T0	vdd	I0/I3081/net13	I0/I3081/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I3058/T0	vdd	I0/I3058/net13	I0/I3058/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2818/T0	vdd	I0/I2818/net13	I0/I2818/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2822/T0	vdd	I0/I2822/net13	I0/I2822/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2817/T0	vdd	I0/I2817/net13	I0/I2817/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2806/T0	vdd	I0/I2806/net13	I0/I2806/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2807/T0	vdd	I0/I2807/net13	I0/I2807/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2818/T1	I0/I2818/net13	I0/I2818/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2822/T1	I0/I2822/net13	I0/I2822/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2817/T1	I0/I2817/net13	I0/I2817/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2806/T1	I0/I2806/net13	I0/I2806/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2807/T1	I0/I2807/net13	I0/I2807/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2870/T0	vdd	I0/I2870/net13	I0/I2870/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2869/T0	vdd	I0/I2869/net13	I0/I2869/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2878/T0	vdd	I0/I2878/net13	I0/I2878/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2884/T0	vdd	I0/I2884/net13	I0/I2884/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2863/T0	vdd	I0/I2863/net13	I0/I2863/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2870/T1	I0/I2870/net13	I0/I2870/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2869/T1	I0/I2869/net13	I0/I2869/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2878/T1	I0/I2878/net13	I0/I2878/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2884/T1	I0/I2884/net13	I0/I2884/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2863/T1	I0/I2863/net13	I0/I2863/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2898/T1	I0/I2898/net13	I0/I2898/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2899/T1	I0/I2899/net13	I0/I2899/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2900/T1	I0/I2900/net13	I0/I2900/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2904/T1	I0/I2904/net13	I0/I2904/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2925/T1	I0/I2925/net13	I0/I2925/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2898/T0	vdd	I0/I2898/net13	I0/I2898/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2899/T0	vdd	I0/I2899/net13	I0/I2899/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2900/T0	vdd	I0/I2900/net13	I0/I2900/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2904/T0	vdd	I0/I2904/net13	I0/I2904/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2925/T0	vdd	I0/I2925/net13	I0/I2925/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2930/T0	vdd	I0/I2930/net13	I0/I2930/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2931/T0	vdd	I0/I2931/net13	I0/I2931/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2927/T0	vdd	I0/I2927/net13	I0/I2927/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2939/T0	vdd	I0/I2939/net13	I0/I2939/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2937/T0	vdd	I0/I2937/net13	I0/I2937/net049	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0504P	AS=0.0896P	PD=0.64U	PS=1.2U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.36e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2930/T1	I0/I2930/net13	I0/I2930/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2931/T1	I0/I2931/net13	I0/I2931/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2927/T1	I0/I2927/net13	I0/I2927/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2939/T1	I0/I2939/net13	I0/I2939/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.24e-14 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.12e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI0/I2937/T1	I0/I2937/net13	I0/I2937/net049	vdd	vdd	pfet
+ L=0.12U	W=0.28U
+ AD=0.0896P	AS=0.0504P	PD=1.2U	PS=0.64U
+ wt=2.8e-07 wf=2.8e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw6=9.6e-15 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=3.36e-14 nrs=0.93617 nrd=0.93617 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI53/T0	BL11	y4bar	net740	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI54/T0	net741	y3bar	BL10bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI55/T0	BL10	y3bar	net740	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI56/T0	net741	y2bar	BL9bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI57/T0	BL9	y2bar	net740	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI58/T0	net741	y1bar	BL8bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI47/T0	BL6	y3bar	net262	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI48/T0	net256	y2bar	BL5bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI49/T0	BL5	y2bar	net262	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI50/T0	net256	y1bar	BL4bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI51/T0	BL4	y1bar	net262	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI52/T0	net741	y4bar	BL11bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI43/T0	net208	y4bar	BL3bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=9.12e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI42/T0	BL3	y4bar	net220	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI41/T0	net208	y3bar	BL2bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI40/T0	BL2	y3bar	net220	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI39/T0	net208	y2bar	BL1bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI38/T0	BL1	y2bar	net220	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI37/T0	net208	y1bar	BL0bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI36/T0	BL0	y1bar	net220	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI44/T0	net256	y4bar	BL7bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI45/T0	BL7	y4bar	net262	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI46/T0	net256	y3bar	BL6bar	vdd	pfet	L=0.12U	W=0.56U
+ AD=0.1792P	AS=0.1792P	PD=1.76U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.6e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=3.6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T3	I116/net60	addr6	vdd	vdd	pfet	L=0.12U
+ W=0.67U
+ AD=0.2144P	AS=0.2144P	PD=1.98U	PS=1.98U
+ wt=6.7e-07 wf=6.7e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.04e-14 panw7=1.044e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.352 nrd=0.352 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T4	I116/net56	I116/net60	vdd	vdd	pfet	L=0.12U
+ W=1.2U
+ AD=0.384P	AS=0.384P	PD=3.04U	PS=3.04U
+ wt=1.2e-06 wf=1.2e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.68e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.2e-14 nrs=0.190476 nrd=0.190476 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T74	y4	I116/net0101	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16U	PS=9.16U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=5.364e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI23/T13	I23/net15	net681	net220	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.64P	PD=2.36U	PS=4.64U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.76e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T12	vdd	I23/net23	I23/net15	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=1.28e-06 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T14	I23/net7	net220	vdd	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.36P	AS=0.36P	PD=2.36U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=8e-07 sa=1.28e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T15	net208	net681	I23/net7	vdd	pfet	L=0.12U
+ W=2U
+ AD=0.64P	AS=0.36P	PD=4.64U	PS=2.36U
+ wt=2e-06 wf=2e-06 sd=0 sb=3.2e-07 sa=1.76e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=2.52e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 panw10=6.6e-14 nrs=0.112532 nrd=0.112532 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T0	vdd	I2/net24	I2/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI2/T1	I2/net20	I2/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI30/T24	I30/net41	I30/net17	vdd	vdd	pfet	L=0.12U
+ W=2.44U
+ AD=0.7808P	AS=0.7808P	PD=5.52U	PS=5.52U
+ wt=2.44e-06 wf=2.44e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.208e-13 nrs=0.091858 nrd=0.091858 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI22/T0	vdd	I22/net24	I22/net24	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=6.72e-14 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T1	I22/net20	I22/net24	vdd	vdd	pfet	L=0.12U
+ W=2.5U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=6.72e-14 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T9	vdd	I22/net20	I22/net8	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1008P	AS=0.1792P	PD=0.92U	PS=1.76U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI22/T10	data0	I22/net8	vdd	vdd	pfet	L=0.12U
+ W=0.56U
+ AD=0.1792P	AS=0.1008P	PD=1.76U	PS=0.92U
+ wt=5.6e-07 wf=5.6e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=7.2e-15 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.427184 nrd=0.427184 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI23/T10	I23/net23	data0	vdd	vdd	pfet	L=0.12U
+ W=0.66U
+ AD=0.2112P	AS=0.2112P	PD=1.96U	PS=1.96U
+ wt=6.6e-07 wf=6.6e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=2.4e-15 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=4.8e-15 nrs=0.357724 nrd=0.357724 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI116/T72	I116/net0101	I116/net0105	vdd	vdd	pfet	L=0.12U
+ W=2.37U
+ AD=0.7584P	AS=0.7584P	PD=5.38U	PS=5.38U
+ wt=2.37e-06 wf=2.37e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=3.072e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0946237 nrd=0.0946237 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T62	vdd	I116/net0281	I116/net0125	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26U	PS=3.26U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.812e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T56	I116/net0281	I116/net120	vdd	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26U	PS=1.17U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.62e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T57	vdd	I116/net0373	I116/net0281	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17U	PS=2.26U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T76	I116/net0229	I116/net0373	vdd	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26U	PS=1.17U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=1.212e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T75	vdd	I116/net56	I116/net0229	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17U	PS=2.26U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.72e-14 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T70	vdd	I116/net0229	I116/net0113	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26U	PS=3.26U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.812e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T71	vdd	I116/net0229	I116/net0105	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26U	PS=3.26U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.461e-13 panw8=5.67e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T73	y4bar	I116/net0113	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16U	PS=9.16U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.352e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T61	vdd	I116/net0281	I116/net0133	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26U	PS=3.26U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.461e-13 panw8=5.67e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T59	y3bar	I116/net0125	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.4058P	PD=9.16U	PS=9.18U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.3e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.352e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T475	vdd	I1/net556	I1/net1744	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T474	I1/net1744	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T464	vdd	I1/net560	I1/net2152	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58U	PS=2.83U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T465	I1/net2152	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83U	PS=5.58U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T476	net929	I1/net1744	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T463	net928	I1/net2152	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.2U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T532	vdd	I1/net1008	I1/net2060	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58001U	PS=2.83001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T531	I1/net2060	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83001U	PS=5.58001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T539	vdd	I1/net1152	I1/net2212	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58001U	PS=2.83001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T540	I1/net2212	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83001U	PS=5.58001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T530	net927	I1/net2060	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.20001U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T538	net926	I1/net2212	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.20001U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T473	I1/net556	I1/net2120	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T466	I1/net560	I1/net1892	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T533	I1/net1008	I1/net2256	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T541	I1/net1152	I1/net2216	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T472	vdd	I1/net1056	I1/net2120	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.40001U	PS=0.74001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T471	I1/net2120	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74001U	PS=0.75001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T470	vdd	I1/a4bar	I1/net2120	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75001U	PS=1.40001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T467	vdd	I1/net1056	I1/net1892	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.40001U	PS=0.74001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T468	I1/net1892	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74001U	PS=0.75001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T469	vdd	I1/a4	I1/net1892	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75001U	PS=1.40001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T536	vdd	I1/net612	I1/net2256	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.40001U	PS=0.74001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T535	I1/net2256	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74001U	PS=0.75001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T534	vdd	I1/a4bar	I1/net2256	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75001U	PS=1.40001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T542	vdd	I1/net612	I1/net2216	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.40001U	PS=0.74001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T543	I1/net2216	I1/a3bar	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74001U	PS=0.75001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T544	vdd	I1/a4	I1/net2216	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75001U	PS=1.40001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T527	vdd	I1/a2	I1/net2184	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.05365P	AS=0.0928P	PD=0.66001U	PS=1.22001U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.03e-14 panw7=2.69e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T528	I1/net2184	I1/a1	vdd	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0522P	AS=0.05365P	PD=0.65001U	PS=0.66001U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=3.48e-14 panw8=8.4e-15 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T537	I1/net612	I1/net2184	vdd	vdd	pfet	L=0.12U
+ W=0.86U
+ AD=0.3096P	AS=0.3182P	PD=2.44001U	PS=2.46001U
+ wt=8.6e-07 wf=8.6e-07 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.224e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.269939 nrd=0.269939 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T529	vdd	I1/a0	I1/net2184	vdd	pfet	L=0.12U
+ W=0.29U
+ AD=0.0928P	AS=0.0522P	PD=1.22001U	PS=0.65001U
+ wt=2.9e-07 wf=2.9e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=4.32e-14 panw7=2.4e-14 panw6=2.4e-15 nrs=0.897959 nrd=0.897959 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=1 PLORIENT=1
MI1/T549	vdd	I1/net612	I1/net2192	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.40001U	PS=0.74001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T550	I1/net2192	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74001U	PS=0.75001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T551	vdd	I1/a4bar	I1/net2192	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75001U	PS=1.40001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T548	I1/net1000	I1/net2192	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T546	vdd	I1/net1000	I1/net2068	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58001U	PS=2.83001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T547	I1/net2068	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83001U	PS=5.58001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T545	net925	I1/net2068	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.20001U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T554	vdd	I1/net612	I1/net2236	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.1216P	AS=0.0684P	PD=1.40001U	PS=0.74001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=3.2e-07 sa=1.29e-06 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=4.56e-14 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T553	I1/net2236	I1/a3	vdd	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0684P	AS=0.0703P	PD=0.74001U	PS=0.75001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=8e-07 sa=8.1e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.56e-14 panw7=9.6e-15 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T552	vdd	I1/a4	I1/net2236	vdd	pfet	L=0.12U
+ W=0.38U
+ AD=0.0703P	AS=0.1216P	PD=0.75001U	PS=1.40001U
+ wt=3.8e-07 wf=3.8e-07 sd=0 sb=1.29e-06 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw7=5.52e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.656716 nrd=0.656716 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T555	I1/net1132	I1/net2236	vdd	vdd	pfet	L=0.12U
+ W=1.12U
+ AD=0.4032P	AS=0.4144P	PD=2.96001U	PS=2.98001U
+ wt=1.12e-06 wf=1.12e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.824e-13 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.4e-15 nrs=0.204651 nrd=0.204651 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T557	vdd	I1/net1132	I1/net2224	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.7904P	AS=0.4446P	PD=5.58001U	PS=2.83001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.74e-14 panw8=2.4e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=3.19e-13 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T556	I1/net2224	I1/addr_en_b	vdd	vdd	pfet	L=0.12U
+ W=2.47U
+ AD=0.4446P	AS=0.7904P	PD=2.83001U	PS=5.58001U
+ wt=2.47e-06 wf=2.47e-06 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.74e-14 panw8=2.71e-13 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=3.6e-15 panw10=7.2e-14 nrs=0.0907216 nrd=0.0907216 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI1/T558	net924	I1/net2224	vdd	vdd	pfet	L=0.12U
+ W=7.24U
+ AD=2.6064P	AS=2.6788P	PD=15.20001U	PS=15.22001U
+ wt=7.24e-06 wf=7.24e-06 sd=0 sb=3.6e-07 sa=3.7e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=5.548e-13 panw8=3.86e-13 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0305768 nrd=0.0305768 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T46	y2	I116/net0145	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16001U	PS=9.16001U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=9.6e-14 panw8=4.8e-14 panw7=5.364e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.44e-13 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T5	I116/net52	addr5	vdd	vdd	pfet	L=0.12U
+ W=0.67U
+ AD=0.2144P	AS=0.2144P	PD=1.98001U	PS=1.98001U
+ wt=6.7e-07 wf=6.7e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.04e-14 panw7=1.044e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.352 nrd=0.352 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T48	I116/net0309	I116/net116	vdd	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26001U	PS=1.17001U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.62e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T6	I116/net0373	I116/net52	vdd	vdd	pfet	L=0.12U
+ W=1.2U
+ AD=0.384P	AS=0.384P	PD=3.04001U	PS=3.04001U
+ wt=1.2e-06 wf=1.2e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.68e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.2e-14 nrs=0.190476 nrd=0.190476 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T0	I116/net120	addr6	vdd	vdd	pfet	L=0.12U
+ W=0.67U
+ AD=0.2144P	AS=0.2144P	PD=1.98001U	PS=1.98001U
+ wt=6.7e-07 wf=6.7e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.04e-14 panw7=1.044e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.352 nrd=0.352 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T14	I116/net96	I116/net116	vdd	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.2592P	AS=0.1458P	PD=2.26001U	PS=1.17001U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=3.2e-07 sa=8e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=1.62e-14 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T1	I116/net116	addr5	vdd	vdd	pfet	L=0.12U
+ W=0.67U
+ AD=0.2144P	AS=0.2144P	PD=1.98001U	PS=1.98001U
+ wt=6.7e-07 wf=6.7e-07 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=2.04e-14 panw7=1.044e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.352 nrd=0.352 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T16	y1	I116/net36	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16001U	PS=9.16001U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.352e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T58	y3	I116/net0137	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16001U	PS=9.16001U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.352e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T44	I116/net0145	I116/net0149	vdd	vdd	pfet	L=0.12U
+ W=2.37U
+ AD=0.7584P	AS=0.7584P	PD=5.38001U	PS=5.38001U
+ wt=2.37e-06 wf=2.37e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=3.072e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0946237 nrd=0.0946237 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T43	vdd	I116/net0309	I116/net0149	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26001U	PS=3.26001U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.461e-13 panw8=5.67e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T45	y2bar	I116/net0157	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16001U	PS=9.16001U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.352e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T42	vdd	I116/net0309	I116/net0157	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26001U	PS=3.26001U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.812e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T47	vdd	I116/net56	I116/net0309	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17001U	PS=2.26001U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T15	vdd	I116/net120	I116/net96	vdd	pfet	L=0.12U
+ W=0.81U
+ AD=0.1458P	AS=0.2592P	PD=1.17001U	PS=2.26001U
+ wt=8.1e-07 wf=8.1e-07 sd=0 sb=8e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw8=3.72e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 nrs=0.287582 nrd=0.287582 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T24	vdd	I116/net96	I116/net24	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26001U	PS=3.26001U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=1.812e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T19	vdd	I116/net96	I116/net32	vdd	pfet	L=0.12U
+ W=1.31U
+ AD=0.4192P	AS=0.4192P	PD=3.26001U	PS=3.26001U
+ wt=1.31e-06 wf=1.31e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=1.461e-13 panw8=5.67e-14 panw7=2.4e-14 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=2.52e-14 nrs=0.173913 nrd=0.173913 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T17	y1bar	I116/net24	vdd	vdd	pfet	L=0.12U
+ W=4.26U
+ AD=1.3632P	AS=1.3632P	PD=9.16001U	PS=9.16001U
+ wt=4.26e-06 wf=4.26e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=5.352e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0521945 nrd=0.0521945 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T18	I116/net36	I116/net32	vdd	vdd	pfet	L=0.12U
+ W=2.37U
+ AD=0.7584P	AS=0.7584P	PD=5.38001U	PS=5.38001U
+ wt=2.37e-06 wf=2.37e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=3.072e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0946237 nrd=0.0946237 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
MI116/T60	I116/net0137	I116/net0133	vdd	vdd	pfet	L=0.12U
+ W=2.37U
+ AD=0.7584P	AS=0.7584P	PD=5.38001U	PS=5.38001U
+ wt=2.37e-06 wf=2.37e-06 sd=0 sb=3.2e-07 sa=3.2e-07 rgatemod=1 rbodymod=0 psp=0 par=1 panw9=4.8e-14 panw8=2.4e-14 panw7=3.072e-13 panw6=1.2e-14 panw5=6e-15 panw4=6e-15 panw3=6e-15 panw2=6e-15 panw10=7.2e-14 nrs=0.0946237 nrd=0.0946237 ngcon=1 nf=1 mSwitch=0 m=1 lstis=1 lnws=1 blockParametersBetween="PC sub" bentgate=0 PWORIENT=0 PLORIENT=0
*
*
*       CAP/DIODE CARDS

*
*       CAPACITOR CARDS
*
*
C1	vdd	vss	1.08059E-12
C2	addr0	vss	7.582E-16
C3	addr1	vss	7.47876E-16
C4	addr2	vss	7.5407E-16
C5	addr3	vss	8.51513E-16
C6	addr4	vss	8.55519E-16
C7	addr5	vss	2.00481E-15
C8	addr6	vss	4.51898E-15
C9	addr_en	vss	4.32417E-16
C10	clk	vss	4.57299E-16
C11	data0	vss	1.16493E-15
C12	data1	vss	1.15315E-15
C13	data2	vss	1.15649E-15
C14	data3	vss	1.15486E-15
C15	data4	vss	1.15764E-15
C16	data5	vss	1.18536E-15
C17	data6	vss	1.18985E-15
C18	data7	vss	1.18703E-15
C19	data8	vss	1.15595E-15
C20	data9	vss	1.15122E-15
C21	wr	vss	1.35861E-15
C22	I1/net148	vss	1.86446E-18
C23	I1/net388	vss	1.75849E-18
C24	I1/net296	vss	1.86446E-18
C25	I1/net584	vss	1.75849E-18
C26	I1/net832	vss	1.86446E-18
C27	I1/net888	vss	1.75849E-18
C28	I1/net840	vss	1.86446E-18
C29	I1/net1048	vss	1.75849E-18
C30	I1/net152	vss	4.54607E-18
C31	I1/net376	vss	4.36154E-18
C32	I1/net512	vss	4.50327E-18
C33	I1/net780	vss	4.34108E-18
C34	I1/net620	vss	4.46083E-18
C35	I1/net884	vss	4.34108E-18
C36	I1/net820	vss	4.46083E-18
C37	I1/net592	vss	4.30042E-18
C38	I1/net168	vss	3.683E-18
C39	I1/net164	vss	4.44828E-18
C40	I1/net108	vss	1.77618E-18
C41	I1/net84	vss	7.04433E-20
C42	I1/net64	vss	1.76841E-18
C43	I1/net380	vss	5.14154E-20
C44	I1/net364	vss	1.77618E-18
C45	I1/net368	vss	7.04433E-20
C46	I1/net340	vss	3.10262E-19
C47	I1/net524	vss	3.683E-18
C48	I1/net520	vss	4.44828E-18
C49	I1/net488	vss	1.77618E-18
C50	I1/net464	vss	7.04433E-20
C51	I1/net444	vss	1.76841E-18
C52	I1/net784	vss	5.14154E-20
C53	I1/net680	vss	1.77618E-18
C54	I1/net692	vss	7.04433E-20
C55	I1/net564	vss	3.10262E-19
C56	I1/net736	vss	3.683E-18
C57	I1/net624	vss	4.44828E-18
C58	I1/net792	vss	1.77618E-18
C59	I1/net660	vss	7.04433E-20
C60	I1/net204	vss	1.76841E-18
C61	I1/net876	vss	5.14154E-20
C62	I1/net912	vss	1.77618E-18
C63	I1/net936	vss	7.04433E-20
C64	I1/net956	vss	3.10262E-19
C65	I1/net1104	vss	3.683E-18
C66	I1/net1060	vss	4.44828E-18
C67	I1/net1124	vss	1.77618E-18
C68	I1/net816	vss	7.04433E-20
C69	I1/net1068	vss	1.76841E-18
C70	I1/net1128	vss	5.14154E-20
C71	I1/net1036	vss	1.77618E-18
C72	I1/net1004	vss	7.04433E-20
C73	I1/net980	vss	3.10262E-19
C74	I1/net984	vss	1.14929E-18
C75	I116/net0326	vss	3.5294E-18
C76	I1/net56	vss	4.59091E-18
C77	I1/net400	vss	4.59091E-18
C78	I1/net436	vss	4.59091E-18
C79	I1/net344	vss	3.54116E-18
C80	I1/net196	vss	4.59091E-18
C81	I1/net964	vss	3.54116E-18
C82	I1/net1080	vss	4.59091E-18
C83	I1/net848	vss	5.43301E-18
C84	I116/net0342	vss	8.52982E-18
C85	I116/net0286	vss	2.91344E-18
C86	I116/net0282	vss	8.48655E-18
C87	I26/net15	vss	1.17844E-15
C88	I0/I3634/net13	vss	7.29973E-16
C89	I0/I3657/net13	vss	7.20083E-16
C90	I0/I4018/net13	vss	7.30111E-16
C91	I0/I3658/net13	vss	7.23918E-16
C92	I0/I4041/net13	vss	7.20083E-16
C93	I0/I3647/net13	vss	7.20083E-16
C94	I0/I4042/net13	vss	7.23918E-16
C95	I0/I3661/net13	vss	7.23918E-16
C96	I0/I4031/net13	vss	7.20083E-16
C97	I0/I3649/net13	vss	7.20083E-16
C98	I0/I4045/net13	vss	7.23918E-16
C99	I0/I3186/net13	vss	7.29973E-16
C100	I0/I3645/net13	vss	7.23918E-16
C101	I0/I4033/net13	vss	7.20083E-16
C102	I0/I3209/net13	vss	7.20083E-16
C103	I0/I3651/net13	vss	7.20083E-16
C104	I0/I4029/net13	vss	7.23918E-16
C105	I0/I3210/net13	vss	7.23918E-16
C106	I0/I3637/net13	vss	7.23918E-16
C107	I0/I4035/net13	vss	7.20083E-16
C108	I0/I3199/net13	vss	7.20083E-16
C109	I0/I3648/net13	vss	7.20083E-16
C110	I0/I4021/net13	vss	7.23918E-16
C111	I0/I3213/net13	vss	7.23918E-16
C112	I0/I3646/net13	vss	7.23918E-16
C113	I0/I4032/net13	vss	7.20083E-16
C114	I0/I3201/net13	vss	7.20083E-16
C115	I0/I3640/net13	vss	7.20083E-16
C116	I0/I4030/net13	vss	7.23918E-16
C117	I0/I3197/net13	vss	7.23918E-16
C118	I0/I3638/net13	vss	7.23918E-16
C119	I0/I4024/net13	vss	7.20083E-16
C120	I0/I3203/net13	vss	7.20083E-16
C121	I0/I3631/net13	vss	7.20083E-16
C122	I0/I4022/net13	vss	7.23918E-16
C123	I0/I3189/net13	vss	7.23918E-16
C124	I0/I3630/net13	vss	7.23918E-16
C125	I0/I4015/net13	vss	7.20083E-16
C126	I0/I3200/net13	vss	7.20083E-16
C127	I0/I3652/net13	vss	7.20083E-16
C128	I0/I4014/net13	vss	7.23918E-16
C129	I0/I3198/net13	vss	7.23918E-16
C130	I0/I3655/net13	vss	7.23918E-16
C131	I0/I4036/net13	vss	7.20083E-16
C132	I0/I3192/net13	vss	7.20083E-16
C133	I0/I3632/net13	vss	7.20083E-16
C134	I0/I4039/net13	vss	7.23918E-16
C135	I0/I3190/net13	vss	7.23918E-16
C136	I0/I3639/net13	vss	7.23918E-16
C137	I0/I4016/net13	vss	7.20083E-16
C138	I0/I3183/net13	vss	7.20083E-16
C139	I0/I3653/net13	vss	7.20083E-16
C140	I0/I4023/net13	vss	7.23918E-16
C141	I0/I3182/net13	vss	7.23918E-16
C142	I0/I3659/net13	vss	7.23918E-16
C143	I0/I4037/net13	vss	7.20083E-16
C144	I0/I3204/net13	vss	7.20083E-16
C145	I0/I3633/net13	vss	7.20083E-16
C146	I0/I4043/net13	vss	7.23918E-16
C147	I0/I3207/net13	vss	7.23918E-16
C148	I0/I3643/net13	vss	7.23918E-16
C149	I0/I4017/net13	vss	7.20083E-16
C150	I0/I3184/net13	vss	7.20083E-16
C151	I0/I3642/net13	vss	7.20083E-16
C152	I0/I4027/net13	vss	7.23918E-16
C153	I0/I3191/net13	vss	7.23918E-16
C154	I0/I3650/net13	vss	7.23918E-16
C155	I0/I4026/net13	vss	7.20083E-16
C156	I0/I3205/net13	vss	7.20083E-16
C157	I0/I3654/net13	vss	7.20083E-16
C158	I0/I4034/net13	vss	7.23918E-16
C159	I0/I3211/net13	vss	7.23918E-16
C160	I0/I3656/net13	vss	7.23918E-16
C161	I0/I4038/net13	vss	7.20083E-16
C162	I0/I3185/net13	vss	7.20083E-16
C163	I0/I3641/net13	vss	7.20083E-16
C164	I0/I4040/net13	vss	7.23918E-16
C165	I0/I3195/net13	vss	7.23918E-16
C166	I0/I3660/net13	vss	7.23918E-16
C167	I0/I4025/net13	vss	7.20083E-16
C168	I0/I3194/net13	vss	7.20083E-16
C169	I0/I3635/net13	vss	7.20083E-16
C170	I0/I4044/net13	vss	7.23918E-16
C171	I0/I3202/net13	vss	7.23918E-16
C172	I0/I3636/net13	vss	7.23918E-16
C173	I0/I4019/net13	vss	7.20083E-16
C174	I0/I3206/net13	vss	7.20083E-16
C175	I0/I3644/net13	vss	7.20313E-16
C176	I0/I4020/net13	vss	7.23918E-16
C177	I0/I3208/net13	vss	7.23918E-16
C178	I0/I4028/net13	vss	7.20313E-16
C179	I0/I3193/net13	vss	7.20083E-16
C180	I0/I3212/net13	vss	7.23918E-16
C181	I0/I3187/net13	vss	7.20083E-16
C182	I0/I3188/net13	vss	7.23918E-16
C183	I0/I3196/net13	vss	7.20313E-16
C184	I22/net8	vss	7.96758E-16
C185	I0/I3634/net049	vss	9.08361E-16
C186	I0/I3657/net049	vss	8.7222E-16
C187	I0/I4018/net049	vss	9.08058E-16
C188	I0/I3658/net049	vss	8.95091E-16
C189	I0/I4041/net049	vss	8.71746E-16
C190	I0/I3647/net049	vss	8.7222E-16
C191	I0/I4042/net049	vss	8.94618E-16
C192	I0/I3661/net049	vss	8.95091E-16
C193	I0/I4031/net049	vss	8.71746E-16
C194	I0/I3649/net049	vss	8.7222E-16
C195	I0/I4045/net049	vss	8.94618E-16
C196	I0/I3186/net049	vss	9.08701E-16
C197	I0/I3645/net049	vss	8.95091E-16
C198	I0/I4033/net049	vss	8.71746E-16
C199	I0/I3209/net049	vss	8.7256E-16
C200	I0/I3651/net049	vss	8.7222E-16
C201	I0/I4029/net049	vss	8.94618E-16
C202	I0/I3210/net049	vss	8.95432E-16
C203	I0/I3637/net049	vss	8.95091E-16
C204	I0/I4035/net049	vss	8.71746E-16
C205	I0/I3199/net049	vss	8.7256E-16
C206	I0/I3648/net049	vss	8.7222E-16
C207	I0/I4021/net049	vss	8.94618E-16
C208	I0/I3213/net049	vss	8.95432E-16
C209	I0/I3646/net049	vss	8.95091E-16
C210	I0/I4032/net049	vss	8.71746E-16
C211	I0/I3201/net049	vss	8.7256E-16
C212	I0/I3640/net049	vss	8.7222E-16
C213	I0/I4030/net049	vss	8.94618E-16
C214	I0/I3197/net049	vss	8.95432E-16
C215	I0/I3638/net049	vss	8.95091E-16
C216	I0/I4024/net049	vss	8.71746E-16
C217	I0/I3203/net049	vss	8.7256E-16
C218	I0/I3631/net049	vss	8.7222E-16
C219	I0/I4022/net049	vss	8.94618E-16
C220	I0/I3189/net049	vss	8.95432E-16
C221	I0/I3630/net049	vss	8.95091E-16
C222	I0/I4015/net049	vss	8.71746E-16
C223	I0/I3200/net049	vss	8.7256E-16
C224	I0/I3652/net049	vss	8.7222E-16
C225	I0/I4014/net049	vss	8.94618E-16
C226	I0/I3198/net049	vss	8.95432E-16
C227	I0/I3655/net049	vss	8.95091E-16
C228	I0/I4036/net049	vss	8.71746E-16
C229	I0/I3192/net049	vss	8.7256E-16
C230	I0/I3632/net049	vss	8.7222E-16
C231	I0/I4039/net049	vss	8.94618E-16
C232	I0/I3190/net049	vss	8.95432E-16
C233	I0/I3639/net049	vss	8.95091E-16
C234	I0/I4016/net049	vss	8.71746E-16
C235	I0/I3183/net049	vss	8.7256E-16
C236	I0/I3653/net049	vss	8.7222E-16
C237	I0/I4023/net049	vss	8.94618E-16
C238	I0/I3182/net049	vss	8.95432E-16
C239	I0/I3659/net049	vss	8.95091E-16
C240	I0/I4037/net049	vss	8.71746E-16
C241	I0/I3204/net049	vss	8.7256E-16
C242	I0/I3633/net049	vss	8.7222E-16
C243	I0/I4043/net049	vss	8.94618E-16
C244	I0/I3207/net049	vss	8.95432E-16
C245	I0/I3643/net049	vss	8.95091E-16
C246	I0/I4017/net049	vss	8.71746E-16
C247	I0/I3184/net049	vss	8.7256E-16
C248	I0/I3642/net049	vss	8.7222E-16
C249	I0/I4027/net049	vss	8.94618E-16
C250	I0/I3191/net049	vss	8.95432E-16
C251	I0/I3650/net049	vss	8.95091E-16
C252	I0/I4026/net049	vss	8.71746E-16
C253	I0/I3205/net049	vss	8.7256E-16
C254	I0/I3654/net049	vss	8.7222E-16
C255	I0/I4034/net049	vss	8.94618E-16
C256	I0/I3211/net049	vss	8.95432E-16
C257	I0/I3656/net049	vss	8.95091E-16
C258	I0/I4038/net049	vss	8.71746E-16
C259	I0/I3185/net049	vss	8.7256E-16
C260	I0/I3641/net049	vss	8.7222E-16
C261	I0/I4040/net049	vss	8.94618E-16
C262	I0/I3195/net049	vss	8.95432E-16
C263	I0/I3660/net049	vss	8.95091E-16
C264	I0/I4025/net049	vss	8.71746E-16
C265	I0/I3194/net049	vss	8.7256E-16
C266	I0/I3635/net049	vss	8.7222E-16
C267	I0/I4044/net049	vss	8.94618E-16
C268	I0/I3202/net049	vss	8.95432E-16
C269	I0/I3636/net049	vss	8.95091E-16
C270	I0/I4019/net049	vss	8.71746E-16
C271	I0/I3206/net049	vss	8.7256E-16
C272	I0/I3644/net049	vss	8.80256E-16
C273	I0/I4020/net049	vss	8.94618E-16
C274	I0/I3208/net049	vss	8.95432E-16
C275	I0/I4028/net049	vss	8.79186E-16
C276	I0/I3193/net049	vss	8.7256E-16
C277	I0/I3212/net049	vss	8.95432E-16
C278	I0/I3187/net049	vss	8.7256E-16
C279	I0/I3188/net049	vss	8.95432E-16
C280	I0/I3196/net049	vss	8.8E-16
C281	I8/net8	vss	7.88667E-16
C282	I22/net20	vss	1.05403E-15
C283	I0/I3410/net13	vss	7.29758E-16
C284	I0/I3433/net13	vss	7.20083E-16
C285	I0/I3794/net13	vss	7.29664E-16
C286	I0/I3434/net13	vss	7.23918E-16
C287	I0/I3817/net13	vss	7.20083E-16
C288	I0/I3423/net13	vss	7.20083E-16
C289	I0/I3818/net13	vss	7.23918E-16
C290	I22/net23	vss	5.28202E-16
C291	I0/I3437/net13	vss	7.23918E-16
C292	I0/I3807/net13	vss	7.20083E-16
C293	I0/I3425/net13	vss	7.20083E-16
C294	I0/I3821/net13	vss	7.23918E-16
C295	I0/I117/net13	vss	7.29758E-16
C296	I0/I3421/net13	vss	7.23918E-16
C297	I0/I3809/net13	vss	7.20083E-16
C298	I0/I94/net13	vss	7.20083E-16
C299	I0/I3427/net13	vss	7.20083E-16
C300	I0/I3805/net13	vss	7.23918E-16
C301	I0/I93/net13	vss	7.23918E-16
C302	I0/I3413/net13	vss	7.23918E-16
C303	I0/I3811/net13	vss	7.20083E-16
C304	I0/I104/net13	vss	7.20083E-16
C305	I0/I3424/net13	vss	7.20083E-16
C306	I0/I3797/net13	vss	7.23918E-16
C307	I0/I90/net13	vss	7.23918E-16
C308	I0/I3422/net13	vss	7.23918E-16
C309	I0/I3808/net13	vss	7.20083E-16
C310	I0/I102/net13	vss	7.20083E-16
C311	I0/I3416/net13	vss	7.20083E-16
C312	I0/I3806/net13	vss	7.23918E-16
C313	I0/I106/net13	vss	7.23918E-16
C314	I0/I3414/net13	vss	7.23918E-16
C315	I0/I3800/net13	vss	7.20083E-16
C316	I0/I100/net13	vss	7.20083E-16
C317	I0/I3407/net13	vss	7.20083E-16
C318	I0/I3798/net13	vss	7.23918E-16
C319	I0/I114/net13	vss	7.23918E-16
C320	I0/I3406/net13	vss	7.23918E-16
C321	I0/I3791/net13	vss	7.20083E-16
C322	I0/I103/net13	vss	7.20083E-16
C323	I0/I3428/net13	vss	7.20083E-16
C324	I0/I3790/net13	vss	7.23918E-16
C325	I0/I105/net13	vss	7.23918E-16
C326	I0/I3431/net13	vss	7.23918E-16
C327	I0/I3812/net13	vss	7.20083E-16
C328	I0/I111/net13	vss	7.20083E-16
C329	I0/I3408/net13	vss	7.20083E-16
C330	I0/I3815/net13	vss	7.23918E-16
C331	I0/I113/net13	vss	7.23918E-16
C332	I0/I3415/net13	vss	7.23918E-16
C333	I0/I3792/net13	vss	7.20083E-16
C334	I0/I120/net13	vss	7.20083E-16
C335	I0/I3429/net13	vss	7.20083E-16
C336	I0/I3799/net13	vss	7.23918E-16
C337	I0/I121/net13	vss	7.23918E-16
C338	I0/I3435/net13	vss	7.23918E-16
C339	I0/I3813/net13	vss	7.20083E-16
C340	I0/I99/net13	vss	7.20083E-16
C341	I0/I3409/net13	vss	7.20083E-16
C342	I0/I3819/net13	vss	7.23918E-16
C343	I0/I96/net13	vss	7.23918E-16
C344	I0/I3419/net13	vss	7.23918E-16
C345	I0/I3793/net13	vss	7.20083E-16
C346	I0/I119/net13	vss	7.20083E-16
C347	I0/I3418/net13	vss	7.20083E-16
C348	I0/I3803/net13	vss	7.23918E-16
C349	I0/I112/net13	vss	7.23918E-16
C350	I0/I3426/net13	vss	7.23918E-16
C351	I0/I3802/net13	vss	7.20083E-16
C352	I0/I98/net13	vss	7.20083E-16
C353	I0/I3430/net13	vss	7.20083E-16
C354	I0/I3810/net13	vss	7.23918E-16
C355	I0/I92/net13	vss	7.23918E-16
C356	I0/I3432/net13	vss	7.23918E-16
C357	I0/I3814/net13	vss	7.20083E-16
C358	I0/I118/net13	vss	7.20083E-16
C359	I0/I3417/net13	vss	7.20083E-16
C360	I0/I3816/net13	vss	7.23918E-16
C361	I0/I108/net13	vss	7.23918E-16
C362	I0/I3436/net13	vss	7.23918E-16
C363	I0/I3801/net13	vss	7.20083E-16
C364	I0/I109/net13	vss	7.20083E-16
C365	I0/I3411/net13	vss	7.20083E-16
C366	I0/I3820/net13	vss	7.23918E-16
C367	I0/I101/net13	vss	7.23918E-16
C368	I0/I3412/net13	vss	7.23918E-16
C369	I0/I3795/net13	vss	7.20083E-16
C370	I0/I97/net13	vss	7.20083E-16
C371	I0/I3420/net13	vss	7.20313E-16
C372	I0/I3796/net13	vss	7.23918E-16
C373	I0/I95/net13	vss	7.23918E-16
C374	I4/net8	vss	7.90771E-16
C375	I0/I3804/net13	vss	7.20313E-16
C376	I0/I110/net13	vss	7.20083E-16
C377	I0/I91/net13	vss	7.23918E-16
C378	I0/I116/net13	vss	7.20083E-16
C379	I0/I115/net13	vss	7.23918E-16
C380	I0/I107/net13	vss	7.20313E-16
C381	I22/net24	vss	6.7709E-16
C382	I0/I3410/net049	vss	9.09062E-16
C383	I8/net20	vss	1.0783E-15
C384	I0/I3433/net049	vss	8.7256E-16
C385	I8/net23	vss	5.26969E-16
C386	I0/I3434/net049	vss	8.95432E-16
C387	I0/I3794/net049	vss	9.08793E-16
C388	I0/I3423/net049	vss	8.7256E-16
C389	I0/I3817/net049	vss	8.7222E-16
C390	I0/I3437/net049	vss	8.95432E-16
C391	I0/I3818/net049	vss	8.95091E-16
C392	I0/I117/net049	vss	9.08578E-16
C393	I0/I3425/net049	vss	8.7256E-16
C394	I0/I3807/net049	vss	8.7222E-16
C395	I0/I94/net049	vss	8.7222E-16
C396	I0/I3421/net049	vss	8.95432E-16
C397	I0/I3821/net049	vss	8.95091E-16
C398	I0/I93/net049	vss	8.95091E-16
C399	I0/I3427/net049	vss	8.7256E-16
C400	I0/I3809/net049	vss	8.7222E-16
C401	I0/I104/net049	vss	8.7222E-16
C402	I0/I3413/net049	vss	8.95432E-16
C403	I0/I3805/net049	vss	8.95091E-16
C404	I0/I90/net049	vss	8.95091E-16
C405	I0/I3424/net049	vss	8.7256E-16
C406	I0/I3811/net049	vss	8.7222E-16
C407	I0/I102/net049	vss	8.7222E-16
C408	I0/I3422/net049	vss	8.95432E-16
C409	I0/I3797/net049	vss	8.95091E-16
C410	I0/I106/net049	vss	8.95091E-16
C411	I0/I3416/net049	vss	8.7256E-16
C412	I0/I3808/net049	vss	8.7222E-16
C413	I0/I100/net049	vss	8.7222E-16
C414	I0/I3414/net049	vss	8.95432E-16
C415	I0/I3806/net049	vss	8.95091E-16
C416	I0/I114/net049	vss	8.95091E-16
C417	I0/I3407/net049	vss	8.7256E-16
C418	I0/I3800/net049	vss	8.7222E-16
C419	I0/I103/net049	vss	8.7222E-16
C420	I0/I3406/net049	vss	8.95432E-16
C421	I0/I3798/net049	vss	8.95091E-16
C422	I0/I105/net049	vss	8.95091E-16
C423	I0/I3428/net049	vss	8.7256E-16
C424	I0/I3791/net049	vss	8.7222E-16
C425	I0/I111/net049	vss	8.7222E-16
C426	I0/I3431/net049	vss	8.95432E-16
C427	I0/I3790/net049	vss	8.95091E-16
C428	I0/I113/net049	vss	8.95091E-16
C429	I0/I3408/net049	vss	8.7256E-16
C430	I0/I3812/net049	vss	8.7222E-16
C431	I0/I120/net049	vss	8.7222E-16
C432	I0/I3415/net049	vss	8.95432E-16
C433	I0/I3815/net049	vss	8.95091E-16
C434	I0/I121/net049	vss	8.95091E-16
C435	I0/I3429/net049	vss	8.7256E-16
C436	I0/I3792/net049	vss	8.7222E-16
C437	I0/I99/net049	vss	8.7222E-16
C438	I0/I3435/net049	vss	8.95432E-16
C439	I0/I3799/net049	vss	8.95091E-16
C440	I0/I96/net049	vss	8.95091E-16
C441	I0/I3409/net049	vss	8.7256E-16
C442	I0/I3813/net049	vss	8.7222E-16
C443	I0/I119/net049	vss	8.7222E-16
C444	I0/I3419/net049	vss	8.95432E-16
C445	I0/I3819/net049	vss	8.95091E-16
C446	I0/I112/net049	vss	8.95091E-16
C447	I0/I3418/net049	vss	8.7256E-16
C448	I0/I3793/net049	vss	8.7222E-16
C449	I0/I98/net049	vss	8.7222E-16
C450	I0/I3426/net049	vss	8.95432E-16
C451	I0/I3803/net049	vss	8.95091E-16
C452	I0/I92/net049	vss	8.95091E-16
C453	I0/I3430/net049	vss	8.7256E-16
C454	I0/I3802/net049	vss	8.7222E-16
C455	I0/I118/net049	vss	8.7222E-16
C456	I0/I3432/net049	vss	8.95432E-16
C457	I0/I3810/net049	vss	8.95091E-16
C458	I0/I108/net049	vss	8.95091E-16
C459	I0/I3417/net049	vss	8.7256E-16
C460	I0/I3814/net049	vss	8.7222E-16
C461	I0/I109/net049	vss	8.7222E-16
C462	I0/I3436/net049	vss	8.95432E-16
C463	I0/I3816/net049	vss	8.95091E-16
C464	I0/I101/net049	vss	8.95091E-16
C465	I0/I3411/net049	vss	8.7256E-16
C466	I0/I3801/net049	vss	8.7222E-16
C467	I0/I97/net049	vss	8.7222E-16
C468	I0/I3412/net049	vss	8.95432E-16
C469	I0/I3820/net049	vss	8.95091E-16
C470	I0/I95/net049	vss	8.95091E-16
C471	I0/I3420/net049	vss	8.8E-16
C472	I0/I3795/net049	vss	8.7222E-16
C473	I0/I110/net049	vss	8.7222E-16
C474	I0/I3796/net049	vss	8.95091E-16
C475	I0/I91/net049	vss	8.95091E-16
C476	I0/I3804/net049	vss	8.79659E-16
C477	I0/I116/net049	vss	8.7222E-16
C478	I0/I115/net049	vss	8.95091E-16
C479	I8/net24	vss	6.8031E-16
C480	I0/I107/net049	vss	8.80256E-16
C481	I4/net20	vss	1.07383E-15
C482	I4/net23	vss	5.34461E-16
C483	I0/I3442/net13	vss	7.29664E-16
C484	I0/I3465/net13	vss	7.20083E-16
C485	I0/I3826/net13	vss	7.29871E-16
C486	I116/net0101	vss	2.54577E-15
C487	I0/I3466/net13	vss	7.23918E-16
C488	I0/I3849/net13	vss	7.20083E-16
C489	I0/I3455/net13	vss	7.20083E-16
C490	I0/I3850/net13	vss	7.23918E-16
C491	I0/I2994/net13	vss	7.29664E-16
C492	I0/I3469/net13	vss	7.23918E-16
C493	I0/I3839/net13	vss	7.20083E-16
C494	I0/I3017/net13	vss	7.20083E-16
C495	I0/I3457/net13	vss	7.20083E-16
C496	I0/I3853/net13	vss	7.23918E-16
C497	I0/I3018/net13	vss	7.23918E-16
C498	I0/I3453/net13	vss	7.23918E-16
C499	I0/I3841/net13	vss	7.20083E-16
C500	I0/I3007/net13	vss	7.20083E-16
C501	I0/I3459/net13	vss	7.20083E-16
C502	I0/I3837/net13	vss	7.23918E-16
C503	I0/I3021/net13	vss	7.23918E-16
C504	I0/I3445/net13	vss	7.23918E-16
C505	I0/I3843/net13	vss	7.20083E-16
C506	I0/I3009/net13	vss	7.20083E-16
C507	I0/I3456/net13	vss	7.20083E-16
C508	I0/I3829/net13	vss	7.23918E-16
C509	I0/I3005/net13	vss	7.23918E-16
C510	I0/I3454/net13	vss	7.23918E-16
C511	I0/I3840/net13	vss	7.20083E-16
C512	I0/I3011/net13	vss	7.20083E-16
C513	I0/I3448/net13	vss	7.20083E-16
C514	I0/I3838/net13	vss	7.23918E-16
C515	I0/I2997/net13	vss	7.23918E-16
C516	I0/I3446/net13	vss	7.23918E-16
C517	I0/I3832/net13	vss	7.20083E-16
C518	I0/I3008/net13	vss	7.20083E-16
C519	I0/I3439/net13	vss	7.20083E-16
C520	I0/I3830/net13	vss	7.23918E-16
C521	I0/I3006/net13	vss	7.23918E-16
C522	I0/I3438/net13	vss	7.23918E-16
C523	I0/I3823/net13	vss	7.20083E-16
C524	I0/I3000/net13	vss	7.20083E-16
C525	I0/I3460/net13	vss	7.20083E-16
C526	I0/I3822/net13	vss	7.23918E-16
C527	I0/I2998/net13	vss	7.23918E-16
C528	I0/I3463/net13	vss	7.23918E-16
C529	I0/I3844/net13	vss	7.20083E-16
C530	I0/I2991/net13	vss	7.20083E-16
C531	I0/I3440/net13	vss	7.20083E-16
C532	I0/I3847/net13	vss	7.23918E-16
C533	I0/I2990/net13	vss	7.23918E-16
C534	I0/I3447/net13	vss	7.23918E-16
C535	I0/I3824/net13	vss	7.20083E-16
C536	I0/I3012/net13	vss	7.20083E-16
C537	I0/I3461/net13	vss	7.20083E-16
C538	I0/I3831/net13	vss	7.23918E-16
C539	I0/I3015/net13	vss	7.23918E-16
C540	I0/I3467/net13	vss	7.23918E-16
C541	I0/I3845/net13	vss	7.20083E-16
C542	I0/I2992/net13	vss	7.20083E-16
C543	I0/I3441/net13	vss	7.20083E-16
C544	I0/I3851/net13	vss	7.23918E-16
C545	I0/I2999/net13	vss	7.23918E-16
C546	I0/I3451/net13	vss	7.23918E-16
C547	I0/I3825/net13	vss	7.20083E-16
C548	I0/I3013/net13	vss	7.20083E-16
C549	I0/I3450/net13	vss	7.20083E-16
C550	I0/I3835/net13	vss	7.23918E-16
C551	I0/I3019/net13	vss	7.23918E-16
C552	I0/I3458/net13	vss	7.23918E-16
C553	I0/I3834/net13	vss	7.20083E-16
C554	I0/I2993/net13	vss	7.20083E-16
C555	I0/I3462/net13	vss	7.20083E-16
C556	I0/I3842/net13	vss	7.23918E-16
C557	I0/I3003/net13	vss	7.23918E-16
C558	I0/I3464/net13	vss	7.23918E-16
C559	I0/I3846/net13	vss	7.20083E-16
C560	I0/I3002/net13	vss	7.20083E-16
C561	I0/I3449/net13	vss	7.20083E-16
C562	I0/I3848/net13	vss	7.23918E-16
C563	I0/I3010/net13	vss	7.23918E-16
C564	I0/I3468/net13	vss	7.23918E-16
C565	I0/I3833/net13	vss	7.20083E-16
C566	I0/I3014/net13	vss	7.20083E-16
C567	I0/I3443/net13	vss	7.20083E-16
C568	I0/I3852/net13	vss	7.23918E-16
C569	I0/I3016/net13	vss	7.23918E-16
C570	I0/I3444/net13	vss	7.23918E-16
C571	I0/I3827/net13	vss	7.20083E-16
C572	I0/I3001/net13	vss	7.20083E-16
C573	I0/I3452/net13	vss	7.20313E-16
C574	I0/I3828/net13	vss	7.23918E-16
C575	I0/I3020/net13	vss	7.23918E-16
C576	I0/I3836/net13	vss	7.20313E-16
C577	I4/net24	vss	6.21617E-16
C578	I0/I2995/net13	vss	7.20083E-16
C579	I29/net7	vss	1.15068E-15
C580	I0/I2996/net13	vss	7.23918E-16
C581	I0/I3004/net13	vss	7.20313E-16
C582	I0/I3442/net049	vss	9.07863E-16
C583	I0/I3465/net049	vss	8.71746E-16
C584	I0/I3826/net049	vss	9.08508E-16
C585	I0/I3466/net049	vss	8.94618E-16
C586	I0/I2994/net049	vss	9.08848E-16
C587	I0/I3849/net049	vss	8.7222E-16
C588	I0/I3455/net049	vss	8.71746E-16
C589	I0/I3017/net049	vss	8.7256E-16
C590	I0/I3469/net049	vss	8.94618E-16
C591	I0/I3850/net049	vss	8.95091E-16
C592	I0/I3018/net049	vss	8.95432E-16
C593	I0/I3457/net049	vss	8.71746E-16
C594	I0/I3839/net049	vss	8.7222E-16
C595	I0/I3007/net049	vss	8.7256E-16
C596	I0/I3453/net049	vss	8.94618E-16
C597	I0/I3853/net049	vss	8.95091E-16
C598	I0/I3021/net049	vss	8.95432E-16
C599	I0/I3459/net049	vss	8.71746E-16
C600	I0/I3841/net049	vss	8.7222E-16
C601	I0/I3009/net049	vss	8.7256E-16
C602	I0/I3445/net049	vss	8.94618E-16
C603	I0/I3837/net049	vss	8.95091E-16
C604	I0/I3005/net049	vss	8.95432E-16
C605	I0/I3456/net049	vss	8.71746E-16
C606	I0/I3843/net049	vss	8.7222E-16
C607	I0/I3011/net049	vss	8.7256E-16
C608	I0/I3454/net049	vss	8.94618E-16
C609	I0/I3829/net049	vss	8.95091E-16
C610	I0/I2997/net049	vss	8.95432E-16
C611	I0/I3448/net049	vss	8.71746E-16
C612	I0/I3840/net049	vss	8.7222E-16
C613	I0/I3008/net049	vss	8.7256E-16
C614	I0/I3446/net049	vss	8.94618E-16
C615	I0/I3838/net049	vss	8.95091E-16
C616	I0/I3006/net049	vss	8.95432E-16
C617	I0/I3439/net049	vss	8.71746E-16
C618	I0/I3832/net049	vss	8.7222E-16
C619	I0/I3000/net049	vss	8.7256E-16
C620	I0/I3438/net049	vss	8.94618E-16
C621	I0/I3830/net049	vss	8.95091E-16
C622	I0/I2998/net049	vss	8.95432E-16
C623	I0/I3460/net049	vss	8.71746E-16
C624	I0/I3823/net049	vss	8.7222E-16
C625	I0/I2991/net049	vss	8.7256E-16
C626	I0/I3463/net049	vss	8.94618E-16
C627	I0/I3822/net049	vss	8.95091E-16
C628	I0/I2990/net049	vss	8.95432E-16
C629	I0/I3440/net049	vss	8.71746E-16
C630	I0/I3844/net049	vss	8.7222E-16
C631	I0/I3012/net049	vss	8.7256E-16
C632	I0/I3447/net049	vss	8.94618E-16
C633	I0/I3847/net049	vss	8.95091E-16
C634	I0/I3015/net049	vss	8.95432E-16
C635	I0/I3461/net049	vss	8.71746E-16
C636	I0/I3824/net049	vss	8.7222E-16
C637	I0/I2992/net049	vss	8.7256E-16
C638	I0/I3467/net049	vss	8.94618E-16
C639	I0/I3831/net049	vss	8.95091E-16
C640	I0/I2999/net049	vss	8.95432E-16
C641	I0/I3441/net049	vss	8.71746E-16
C642	I0/I3845/net049	vss	8.7222E-16
C643	I0/I3013/net049	vss	8.7256E-16
C644	I0/I3451/net049	vss	8.94618E-16
C645	I0/I3851/net049	vss	8.95091E-16
C646	I0/I3019/net049	vss	8.95432E-16
C647	I0/I3450/net049	vss	8.71746E-16
C648	I0/I3825/net049	vss	8.7222E-16
C649	I0/I2993/net049	vss	8.7256E-16
C650	I0/I3458/net049	vss	8.94618E-16
C651	I0/I3835/net049	vss	8.95091E-16
C652	I0/I3003/net049	vss	8.95432E-16
C653	I0/I3462/net049	vss	8.71746E-16
C654	I0/I3834/net049	vss	8.7222E-16
C655	I0/I3002/net049	vss	8.7256E-16
C656	I0/I3464/net049	vss	8.94618E-16
C657	I0/I3842/net049	vss	8.95091E-16
C658	I0/I3010/net049	vss	8.95432E-16
C659	I0/I3449/net049	vss	8.71746E-16
C660	I0/I3846/net049	vss	8.7222E-16
C661	I0/I3014/net049	vss	8.7256E-16
C662	I0/I3468/net049	vss	8.94618E-16
C663	I0/I3848/net049	vss	8.95091E-16
C664	I0/I3016/net049	vss	8.95432E-16
C665	I0/I3443/net049	vss	8.71746E-16
C666	I0/I3833/net049	vss	8.7222E-16
C667	I0/I3001/net049	vss	8.7256E-16
C668	I0/I3444/net049	vss	8.94618E-16
C669	I0/I3852/net049	vss	8.95091E-16
C670	I0/I3020/net049	vss	8.95432E-16
C671	I0/I3452/net049	vss	8.79186E-16
C672	I0/I3827/net049	vss	8.7222E-16
C673	I0/I2995/net049	vss	8.7256E-16
C674	I0/I3828/net049	vss	8.95091E-16
C675	I0/I2996/net049	vss	8.95432E-16
C676	I0/I3836/net049	vss	8.79659E-16
C677	I0/I3004/net049	vss	8.80596E-16
C678	I29/net15	vss	1.18751E-15
C679	I0/I3474/net13	vss	7.29699E-16
C680	I0/I3497/net13	vss	7.20083E-16
C681	I0/I3498/net13	vss	7.23918E-16
C682	I0/I3026/net13	vss	7.29837E-16
C683	I0/I3858/net13	vss	7.29837E-16
C684	I0/I3487/net13	vss	7.20083E-16
C685	I0/I3049/net13	vss	7.20083E-16
C686	I0/I3501/net13	vss	7.23918E-16
C687	I0/I3881/net13	vss	7.20083E-16
C688	I0/I3050/net13	vss	7.23918E-16
C689	I0/I3489/net13	vss	7.20083E-16
C690	I0/I3882/net13	vss	7.23918E-16
C691	I0/I3039/net13	vss	7.20083E-16
C692	I0/I3485/net13	vss	7.23918E-16
C693	I0/I3871/net13	vss	7.20083E-16
C694	I0/I3053/net13	vss	7.23918E-16
C695	I0/I3491/net13	vss	7.20083E-16
C696	I0/I3885/net13	vss	7.23918E-16
C697	I0/I3041/net13	vss	7.20083E-16
C698	I0/I3477/net13	vss	7.23918E-16
C699	I0/I3873/net13	vss	7.20083E-16
C700	I0/I3037/net13	vss	7.23918E-16
C701	I0/I3488/net13	vss	7.20083E-16
C702	I0/I3869/net13	vss	7.23918E-16
C703	I0/I3043/net13	vss	7.20083E-16
C704	I0/I3486/net13	vss	7.23918E-16
C705	I0/I3875/net13	vss	7.20083E-16
C706	I0/I3029/net13	vss	7.23918E-16
C707	I0/I3480/net13	vss	7.20083E-16
C708	I0/I3861/net13	vss	7.23918E-16
C709	I0/I3040/net13	vss	7.20083E-16
C710	I0/I3478/net13	vss	7.23918E-16
C711	I0/I3872/net13	vss	7.20083E-16
C712	I0/I3038/net13	vss	7.23918E-16
C713	I0/I3471/net13	vss	7.20083E-16
C714	I0/I3870/net13	vss	7.23918E-16
C715	I0/I3032/net13	vss	7.20083E-16
C716	I0/I3470/net13	vss	7.23918E-16
C717	I0/I3864/net13	vss	7.20083E-16
C718	I0/I3030/net13	vss	7.23918E-16
C719	I0/I3492/net13	vss	7.20083E-16
C720	I0/I3862/net13	vss	7.23918E-16
C721	I0/I3023/net13	vss	7.20083E-16
C722	I0/I3495/net13	vss	7.23918E-16
C723	I0/I3855/net13	vss	7.20083E-16
C724	I0/I3022/net13	vss	7.23918E-16
C725	I0/I3472/net13	vss	7.20083E-16
C726	I0/I3854/net13	vss	7.23918E-16
C727	I0/I3044/net13	vss	7.20083E-16
C728	I0/I3479/net13	vss	7.23918E-16
C729	I0/I3876/net13	vss	7.20083E-16
C730	I0/I3047/net13	vss	7.23918E-16
C731	I0/I3493/net13	vss	7.20083E-16
C732	I0/I3879/net13	vss	7.23918E-16
C733	I0/I3024/net13	vss	7.20083E-16
C734	I0/I3499/net13	vss	7.23918E-16
C735	I0/I3856/net13	vss	7.20083E-16
C736	I0/I3031/net13	vss	7.23918E-16
C737	I0/I3473/net13	vss	7.20083E-16
C738	I0/I3863/net13	vss	7.23918E-16
C739	I0/I3045/net13	vss	7.20083E-16
C740	I0/I3483/net13	vss	7.23918E-16
C741	I0/I3877/net13	vss	7.20083E-16
C742	I0/I3051/net13	vss	7.23918E-16
C743	I0/I3482/net13	vss	7.20083E-16
C744	I0/I3883/net13	vss	7.23918E-16
C745	I0/I3025/net13	vss	7.20083E-16
C746	I0/I3490/net13	vss	7.23918E-16
C747	I0/I3857/net13	vss	7.20083E-16
C748	I0/I3035/net13	vss	7.23918E-16
C749	I0/I3494/net13	vss	7.20083E-16
C750	I0/I3867/net13	vss	7.23918E-16
C751	I0/I3034/net13	vss	7.20083E-16
C752	I0/I3496/net13	vss	7.23918E-16
C753	I0/I3866/net13	vss	7.20083E-16
C754	I0/I3042/net13	vss	7.23918E-16
C755	I0/I3481/net13	vss	7.20083E-16
C756	I0/I3874/net13	vss	7.23918E-16
C757	I0/I3046/net13	vss	7.20083E-16
C758	I0/I3500/net13	vss	7.23918E-16
C759	I0/I3878/net13	vss	7.20083E-16
C760	I0/I3048/net13	vss	7.23918E-16
C761	I0/I3475/net13	vss	7.20083E-16
C762	I0/I3880/net13	vss	7.23918E-16
C763	I0/I3033/net13	vss	7.20083E-16
C764	I0/I3476/net13	vss	7.23918E-16
C765	I0/I3865/net13	vss	7.20083E-16
C766	I0/I3052/net13	vss	7.23918E-16
C767	I0/I3484/net13	vss	7.20313E-16
C768	I0/I3884/net13	vss	7.23918E-16
C769	I0/I3027/net13	vss	7.20083E-16
C770	I0/I3859/net13	vss	7.20083E-16
C771	I0/I3028/net13	vss	7.23918E-16
C772	I0/I3860/net13	vss	7.23918E-16
C773	I0/I3036/net13	vss	7.20313E-16
C774	I0/I3868/net13	vss	7.20313E-16
C775	I0/I3474/net049	vss	9.09518E-16
C776	I0/I3497/net049	vss	8.71746E-16
C777	I0/I3498/net049	vss	8.94618E-16
C778	I0/I3026/net049	vss	9.09689E-16
C779	I0/I3487/net049	vss	8.71746E-16
C780	I0/I3049/net049	vss	8.71746E-16
C781	I0/I3501/net049	vss	8.94618E-16
C782	I0/I3050/net049	vss	8.94618E-16
C783	I0/I3489/net049	vss	8.71746E-16
C784	I0/I3858/net049	vss	9.09689E-16
C785	I0/I3039/net049	vss	8.71746E-16
C786	I0/I3485/net049	vss	8.94618E-16
C787	I0/I3881/net049	vss	8.71746E-16
C788	I0/I3053/net049	vss	8.94618E-16
C789	I0/I3491/net049	vss	8.71746E-16
C790	I0/I3882/net049	vss	8.94618E-16
C791	I0/I3041/net049	vss	8.71746E-16
C792	I0/I3477/net049	vss	8.94618E-16
C793	I0/I3871/net049	vss	8.71746E-16
C794	I0/I3037/net049	vss	8.94618E-16
C795	I0/I3488/net049	vss	8.71746E-16
C796	I0/I3885/net049	vss	8.94618E-16
C797	I0/I3043/net049	vss	8.71746E-16
C798	I0/I3486/net049	vss	8.94618E-16
C799	I0/I3873/net049	vss	8.71746E-16
C800	I0/I3029/net049	vss	8.94618E-16
C801	I0/I3480/net049	vss	8.71746E-16
C802	I0/I3869/net049	vss	8.94618E-16
C803	I0/I3040/net049	vss	8.71746E-16
C804	I0/I3478/net049	vss	8.94618E-16
C805	I0/I3875/net049	vss	8.71746E-16
C806	I0/I3038/net049	vss	8.94618E-16
C807	I0/I3471/net049	vss	8.71746E-16
C808	I0/I3861/net049	vss	8.94618E-16
C809	I0/I3032/net049	vss	8.71746E-16
C810	I0/I3470/net049	vss	8.94618E-16
C811	I0/I3872/net049	vss	8.71746E-16
C812	I0/I3030/net049	vss	8.94618E-16
C813	I0/I3492/net049	vss	8.71746E-16
C814	I0/I3870/net049	vss	8.94618E-16
C815	I0/I3023/net049	vss	8.71746E-16
C816	I0/I3495/net049	vss	8.94618E-16
C817	I0/I3864/net049	vss	8.71746E-16
C818	I0/I3022/net049	vss	8.94618E-16
C819	I0/I3472/net049	vss	8.71746E-16
C820	I0/I3862/net049	vss	8.94618E-16
C821	I0/I3044/net049	vss	8.71746E-16
C822	I0/I3479/net049	vss	8.94618E-16
C823	I0/I3855/net049	vss	8.71746E-16
C824	I0/I3047/net049	vss	8.94618E-16
C825	I0/I3493/net049	vss	8.71746E-16
C826	I0/I3854/net049	vss	8.94618E-16
C827	I0/I3024/net049	vss	8.71746E-16
C828	I0/I3499/net049	vss	8.94618E-16
C829	I0/I3876/net049	vss	8.71746E-16
C830	I0/I3031/net049	vss	8.94618E-16
C831	I0/I3473/net049	vss	8.71746E-16
C832	I0/I3879/net049	vss	8.94618E-16
C833	I0/I3045/net049	vss	8.71746E-16
C834	I0/I3483/net049	vss	8.94618E-16
C835	I0/I3856/net049	vss	8.71746E-16
C836	I0/I3051/net049	vss	8.94618E-16
C837	I0/I3482/net049	vss	8.71746E-16
C838	I0/I3863/net049	vss	8.94618E-16
C839	I0/I3025/net049	vss	8.71746E-16
C840	I0/I3490/net049	vss	8.94618E-16
C841	I0/I3877/net049	vss	8.71746E-16
C842	I0/I3035/net049	vss	8.94618E-16
C843	I0/I3494/net049	vss	8.71746E-16
C844	I0/I3883/net049	vss	8.94618E-16
C845	I0/I3034/net049	vss	8.71746E-16
C846	I0/I3496/net049	vss	8.94618E-16
C847	I0/I3857/net049	vss	8.71746E-16
C848	I0/I3042/net049	vss	8.94618E-16
C849	I0/I3481/net049	vss	8.71746E-16
C850	I0/I3867/net049	vss	8.94618E-16
C851	I0/I3046/net049	vss	8.71746E-16
C852	I0/I3500/net049	vss	8.94618E-16
C853	I0/I3866/net049	vss	8.71746E-16
C854	I0/I3048/net049	vss	8.94618E-16
C855	I0/I3475/net049	vss	8.71746E-16
C856	I0/I3874/net049	vss	8.94618E-16
C857	I0/I3033/net049	vss	8.71746E-16
C858	I0/I3476/net049	vss	8.94618E-16
C859	I0/I3878/net049	vss	8.71746E-16
C860	I0/I3052/net049	vss	8.94618E-16
C861	I0/I3484/net049	vss	8.79783E-16
C862	I0/I3880/net049	vss	8.94618E-16
C863	I0/I3027/net049	vss	8.71746E-16
C864	I0/I3865/net049	vss	8.71746E-16
C865	I0/I3028/net049	vss	8.94618E-16
C866	I0/I3884/net049	vss	8.94618E-16
C867	I0/I3036/net049	vss	8.79783E-16
C868	I0/I3859/net049	vss	8.71746E-16
C869	I0/I3860/net049	vss	8.94618E-16
C870	I0/I3868/net049	vss	8.79186E-16
C871	I7/net8	vss	7.86207E-16
C872	I25/net7	vss	1.15705E-15
C873	I0/I3506/net13	vss	7.29973E-16
C874	I0/I3058/net13	vss	7.30111E-16
C875	I0/I3529/net13	vss	7.20083E-16
C876	I0/I3081/net13	vss	7.20083E-16
C877	I0/I3530/net13	vss	7.23918E-16
C878	I0/I3082/net13	vss	7.23918E-16
C879	I0/I3519/net13	vss	7.20083E-16
C880	I0/I3071/net13	vss	7.20083E-16
C881	I0/I3533/net13	vss	7.23918E-16
C882	I0/I3085/net13	vss	7.23918E-16
C883	I0/I3521/net13	vss	7.20083E-16
C884	I0/I3073/net13	vss	7.20083E-16
C885	I0/I3517/net13	vss	7.23918E-16
C886	I0/I3069/net13	vss	7.23918E-16
C887	I0/I3523/net13	vss	7.20083E-16
C888	I0/I3890/net13	vss	7.30111E-16
C889	I0/I3075/net13	vss	7.20083E-16
C890	I0/I3509/net13	vss	7.23918E-16
C891	I0/I3913/net13	vss	7.20083E-16
C892	I0/I3061/net13	vss	7.23918E-16
C893	I0/I3520/net13	vss	7.20083E-16
C894	I0/I3914/net13	vss	7.23918E-16
C895	I0/I3072/net13	vss	7.20083E-16
C896	I0/I3518/net13	vss	7.23918E-16
C897	I0/I3903/net13	vss	7.20083E-16
C898	I0/I3070/net13	vss	7.23918E-16
C899	I0/I3512/net13	vss	7.20083E-16
C900	I0/I3917/net13	vss	7.23918E-16
C901	I0/I3064/net13	vss	7.20083E-16
C902	I0/I3510/net13	vss	7.23918E-16
C903	I0/I3905/net13	vss	7.20083E-16
C904	I0/I3062/net13	vss	7.23918E-16
C905	I0/I3503/net13	vss	7.20083E-16
C906	I0/I3901/net13	vss	7.23918E-16
C907	I0/I3055/net13	vss	7.20083E-16
C908	I0/I3502/net13	vss	7.23918E-16
C909	I0/I3907/net13	vss	7.20083E-16
C910	I0/I3054/net13	vss	7.23918E-16
C911	I0/I3524/net13	vss	7.20083E-16
C912	I0/I3893/net13	vss	7.23918E-16
C913	I0/I3076/net13	vss	7.20083E-16
C914	I0/I3527/net13	vss	7.23918E-16
C915	I0/I3904/net13	vss	7.20083E-16
C916	I0/I3079/net13	vss	7.23918E-16
C917	I0/I3504/net13	vss	7.20083E-16
C918	I0/I3902/net13	vss	7.23918E-16
C919	I0/I3056/net13	vss	7.20083E-16
C920	I0/I3511/net13	vss	7.23918E-16
C921	I0/I3896/net13	vss	7.20083E-16
C922	I0/I3063/net13	vss	7.23918E-16
C923	I0/I3525/net13	vss	7.20083E-16
C924	I0/I3894/net13	vss	7.23918E-16
C925	I0/I3077/net13	vss	7.20083E-16
C926	I0/I3531/net13	vss	7.23918E-16
C927	I0/I3887/net13	vss	7.20083E-16
C928	I0/I3083/net13	vss	7.23918E-16
C929	I0/I3505/net13	vss	7.20083E-16
C930	I0/I3886/net13	vss	7.23918E-16
C931	I0/I3057/net13	vss	7.20083E-16
C932	I0/I3515/net13	vss	7.23918E-16
C933	I0/I3908/net13	vss	7.20083E-16
C934	I0/I3067/net13	vss	7.23918E-16
C935	I0/I3514/net13	vss	7.20083E-16
C936	I0/I3911/net13	vss	7.23918E-16
C937	I0/I3066/net13	vss	7.20083E-16
C938	I0/I3522/net13	vss	7.23918E-16
C939	I0/I3888/net13	vss	7.20083E-16
C940	I0/I3074/net13	vss	7.23918E-16
C941	I0/I3526/net13	vss	7.20083E-16
C942	I0/I3895/net13	vss	7.23918E-16
C943	I0/I3078/net13	vss	7.20083E-16
C944	I0/I3528/net13	vss	7.23918E-16
C945	I0/I3909/net13	vss	7.20083E-16
C946	I0/I3080/net13	vss	7.23918E-16
C947	I0/I3513/net13	vss	7.20083E-16
C948	I0/I3915/net13	vss	7.23918E-16
C949	I0/I3065/net13	vss	7.20083E-16
C950	I0/I3532/net13	vss	7.23918E-16
C951	I0/I3889/net13	vss	7.20083E-16
C952	I0/I3084/net13	vss	7.23918E-16
C953	I0/I3507/net13	vss	7.20083E-16
C954	I0/I3899/net13	vss	7.23918E-16
C955	I0/I3059/net13	vss	7.20083E-16
C956	I0/I3508/net13	vss	7.23918E-16
C957	I0/I3898/net13	vss	7.20083E-16
C958	I0/I3060/net13	vss	7.23918E-16
C959	I0/I3516/net13	vss	7.20313E-16
C960	I0/I3906/net13	vss	7.23918E-16
C961	I0/I3068/net13	vss	7.20313E-16
C962	I0/I3910/net13	vss	7.20083E-16
C963	I0/I3912/net13	vss	7.23918E-16
C964	I0/I3897/net13	vss	7.20083E-16
C965	I0/I3916/net13	vss	7.23918E-16
C966	I0/I3891/net13	vss	7.20083E-16
C967	I0/I3892/net13	vss	7.23918E-16
C968	I0/I3900/net13	vss	7.20313E-16
C969	I25/net15	vss	1.17512E-15
C970	I0/I3506/net049	vss	9.08701E-16
C971	I0/I3058/net049	vss	9.08872E-16
C972	I0/I3529/net049	vss	8.7256E-16
C973	I0/I3081/net049	vss	8.7256E-16
C974	I0/I3530/net049	vss	8.95432E-16
C975	I0/I3082/net049	vss	8.95432E-16
C976	I0/I3519/net049	vss	8.7256E-16
C977	I0/I3071/net049	vss	8.7256E-16
C978	I0/I3533/net049	vss	8.95432E-16
C979	I0/I3085/net049	vss	8.95432E-16
C980	I7/net20	vss	1.07497E-15
C981	I0/I3521/net049	vss	8.7256E-16
C982	I0/I3073/net049	vss	8.7256E-16
C983	I7/net23	vss	5.32741E-16
C984	I0/I3517/net049	vss	8.95432E-16
C985	I0/I3069/net049	vss	8.95432E-16
C986	I0/I3890/net049	vss	9.08787E-16
C987	I0/I3523/net049	vss	8.7256E-16
C988	I0/I3075/net049	vss	8.7256E-16
C989	I0/I3913/net049	vss	8.7256E-16
C990	I0/I3509/net049	vss	8.95432E-16
C991	I0/I3061/net049	vss	8.95432E-16
C992	I0/I3914/net049	vss	8.95432E-16
C993	I0/I3520/net049	vss	8.7256E-16
C994	I0/I3072/net049	vss	8.7256E-16
C995	I0/I3903/net049	vss	8.7256E-16
C996	I0/I3518/net049	vss	8.95432E-16
C997	I0/I3070/net049	vss	8.95432E-16
C998	I0/I3917/net049	vss	8.95432E-16
C999	I0/I3512/net049	vss	8.7256E-16
C1000	I0/I3064/net049	vss	8.7256E-16
C1001	I0/I3510/net049	vss	8.95432E-16
C1002	I0/I3905/net049	vss	8.7256E-16
C1003	I0/I3062/net049	vss	8.95432E-16
C1004	I0/I3503/net049	vss	8.7256E-16
C1005	I0/I3901/net049	vss	8.95432E-16
C1006	I0/I3055/net049	vss	8.7256E-16
C1007	I0/I3502/net049	vss	8.95432E-16
C1008	I0/I3907/net049	vss	8.7256E-16
C1009	I0/I3054/net049	vss	8.95432E-16
C1010	I0/I3524/net049	vss	8.7256E-16
C1011	I0/I3893/net049	vss	8.95432E-16
C1012	I0/I3076/net049	vss	8.7256E-16
C1013	I0/I3527/net049	vss	8.95432E-16
C1014	I0/I3904/net049	vss	8.7256E-16
C1015	I0/I3079/net049	vss	8.95432E-16
C1016	I0/I3504/net049	vss	8.7256E-16
C1017	I0/I3902/net049	vss	8.95432E-16
C1018	I0/I3056/net049	vss	8.7256E-16
C1019	I0/I3511/net049	vss	8.95432E-16
C1020	I0/I3896/net049	vss	8.7256E-16
C1021	I0/I3063/net049	vss	8.95432E-16
C1022	I0/I3525/net049	vss	8.7256E-16
C1023	I0/I3894/net049	vss	8.95432E-16
C1024	I0/I3077/net049	vss	8.7256E-16
C1025	I0/I3531/net049	vss	8.95432E-16
C1026	I0/I3887/net049	vss	8.7256E-16
C1027	I0/I3083/net049	vss	8.95432E-16
C1028	I0/I3505/net049	vss	8.7256E-16
C1029	I0/I3886/net049	vss	8.95432E-16
C1030	I0/I3057/net049	vss	8.7256E-16
C1031	I0/I3515/net049	vss	8.95432E-16
C1032	I0/I3908/net049	vss	8.7256E-16
C1033	I0/I3067/net049	vss	8.95432E-16
C1034	I0/I3514/net049	vss	8.7256E-16
C1035	I0/I3911/net049	vss	8.95432E-16
C1036	I0/I3066/net049	vss	8.7256E-16
C1037	I0/I3522/net049	vss	8.95432E-16
C1038	I0/I3888/net049	vss	8.7256E-16
C1039	I0/I3074/net049	vss	8.95432E-16
C1040	I0/I3526/net049	vss	8.7256E-16
C1041	I0/I3895/net049	vss	8.95432E-16
C1042	I0/I3078/net049	vss	8.7256E-16
C1043	I0/I3528/net049	vss	8.95432E-16
C1044	I0/I3909/net049	vss	8.7256E-16
C1045	I0/I3080/net049	vss	8.95432E-16
C1046	I0/I3513/net049	vss	8.7256E-16
C1047	I0/I3915/net049	vss	8.95432E-16
C1048	I0/I3065/net049	vss	8.7256E-16
C1049	I0/I3532/net049	vss	8.95432E-16
C1050	I0/I3889/net049	vss	8.7256E-16
C1051	I0/I3084/net049	vss	8.95432E-16
C1052	I0/I3507/net049	vss	8.7256E-16
C1053	I0/I3899/net049	vss	8.95432E-16
C1054	I0/I3059/net049	vss	8.7256E-16
C1055	I0/I3508/net049	vss	8.95432E-16
C1056	I0/I3898/net049	vss	8.7256E-16
C1057	I0/I3060/net049	vss	8.95432E-16
C1058	I0/I3516/net049	vss	8.80596E-16
C1059	I0/I3906/net049	vss	8.95432E-16
C1060	I0/I3068/net049	vss	8.80596E-16
C1061	I0/I3910/net049	vss	8.7256E-16
C1062	I0/I3912/net049	vss	8.95432E-16
C1063	I0/I3897/net049	vss	8.7256E-16
C1064	I0/I3916/net049	vss	8.95432E-16
C1065	I0/I3891/net049	vss	8.7256E-16
C1066	I0/I3892/net049	vss	8.95432E-16
C1067	I0/I3900/net049	vss	8.8E-16
C1068	I7/net24	vss	6.83342E-16
C1069	I116/net0105	vss	2.09176E-15
C1070	I0/I2807/net13	vss	7.29871E-16
C1071	I0/I2806/net13	vss	7.20083E-16
C1072	I0/I2817/net13	vss	7.23918E-16
C1073	I0/I3282/net13	vss	7.29758E-16
C1074	I0/I2822/net13	vss	7.20083E-16
C1075	I0/I3305/net13	vss	7.20083E-16
C1076	I0/I2818/net13	vss	7.23918E-16
C1077	I0/I3306/net13	vss	7.23918E-16
C1078	I0/I2814/net13	vss	7.20083E-16
C1079	I0/I4050/net13	vss	7.42504E-16
C1080	I0/I3295/net13	vss	7.20083E-16
C1081	I0/I2815/net13	vss	7.23918E-16
C1082	I0/I3666/net13	vss	7.29656E-16
C1083	I0/I4073/net13	vss	7.44139E-16
C1084	I0/I3309/net13	vss	7.23918E-16
C1085	I0/I2819/net13	vss	7.20083E-16
C1086	I0/I3689/net13	vss	7.20083E-16
C1087	I0/I4074/net13	vss	7.42366E-16
C1088	I0/I3297/net13	vss	7.20083E-16
C1089	I0/I2808/net13	vss	7.23918E-16
C1090	I0/I3690/net13	vss	7.23918E-16
C1091	I0/I4063/net13	vss	7.44139E-16
C1092	I0/I3293/net13	vss	7.23918E-16
C1093	I0/I2824/net13	vss	7.20083E-16
C1094	I0/I3679/net13	vss	7.20083E-16
C1095	I0/I4077/net13	vss	7.42366E-16
C1096	I0/I3299/net13	vss	7.20083E-16
C1097	I0/I2823/net13	vss	7.23918E-16
C1098	I0/I3693/net13	vss	7.23918E-16
C1099	I0/I4065/net13	vss	7.44139E-16
C1100	I0/I3285/net13	vss	7.23918E-16
C1101	I0/I2801/net13	vss	7.20083E-16
C1102	I0/I3681/net13	vss	7.20083E-16
C1103	I0/I4061/net13	vss	7.42366E-16
C1104	I0/I3296/net13	vss	7.20083E-16
C1105	I0/I2809/net13	vss	7.23918E-16
C1106	I0/I3677/net13	vss	7.23918E-16
C1107	I0/I4067/net13	vss	7.44139E-16
C1108	I0/I3294/net13	vss	7.23918E-16
C1109	I0/I2810/net13	vss	7.20083E-16
C1110	I0/I3683/net13	vss	7.20083E-16
C1111	I0/I4053/net13	vss	7.42366E-16
C1112	I0/I3288/net13	vss	7.20083E-16
C1113	I0/I2800/net13	vss	7.23918E-16
C1114	I0/I3669/net13	vss	7.23918E-16
C1115	I0/I4064/net13	vss	7.44139E-16
C1116	I0/I3286/net13	vss	7.23918E-16
C1117	I0/I2820/net13	vss	7.20083E-16
C1118	I0/I3279/net13	vss	7.20083E-16
C1119	I0/I3680/net13	vss	7.20083E-16
C1120	I0/I4062/net13	vss	7.42366E-16
C1121	I0/I2802/net13	vss	7.23918E-16
C1122	I0/I3278/net13	vss	7.23918E-16
C1123	I0/I3678/net13	vss	7.23918E-16
C1124	I0/I4056/net13	vss	7.44139E-16
C1125	I0/I2804/net13	vss	7.20083E-16
C1126	I0/I3300/net13	vss	7.20083E-16
C1127	I0/I3672/net13	vss	7.20083E-16
C1128	I0/I4054/net13	vss	7.42366E-16
C1129	I0/I2827/net13	vss	7.23918E-16
C1130	I0/I3303/net13	vss	7.23918E-16
C1131	I0/I3670/net13	vss	7.23918E-16
C1132	I0/I4047/net13	vss	7.44139E-16
C1133	I0/I2813/net13	vss	7.20083E-16
C1134	I0/I3280/net13	vss	7.20083E-16
C1135	I0/I3663/net13	vss	7.20083E-16
C1136	I0/I4046/net13	vss	7.42366E-16
C1137	I0/I2811/net13	vss	7.23918E-16
C1138	I0/I3287/net13	vss	7.23918E-16
C1139	I0/I3662/net13	vss	7.23918E-16
C1140	I0/I4068/net13	vss	7.44139E-16
C1141	I0/I2803/net13	vss	7.20083E-16
C1142	I0/I3301/net13	vss	7.20083E-16
C1143	I0/I3684/net13	vss	7.20083E-16
C1144	I0/I4071/net13	vss	7.42366E-16
C1145	I0/I2816/net13	vss	7.23918E-16
C1146	I0/I3307/net13	vss	7.23918E-16
C1147	I0/I3687/net13	vss	7.23918E-16
C1148	I0/I4048/net13	vss	7.44139E-16
C1149	I0/I2826/net13	vss	7.20083E-16
C1150	I0/I3281/net13	vss	7.20083E-16
C1151	I0/I3664/net13	vss	7.20083E-16
C1152	I0/I4055/net13	vss	7.42366E-16
C1153	I0/I2805/net13	vss	7.23918E-16
C1154	I0/I3291/net13	vss	7.23918E-16
C1155	I0/I3671/net13	vss	7.23918E-16
C1156	I0/I4069/net13	vss	7.44139E-16
C1157	I0/I2825/net13	vss	7.20083E-16
C1158	I0/I3290/net13	vss	7.20083E-16
C1159	I0/I3685/net13	vss	7.20083E-16
C1160	I0/I4075/net13	vss	7.42366E-16
C1161	I0/I2812/net13	vss	7.23918E-16
C1162	I0/I3298/net13	vss	7.23918E-16
C1163	I0/I3691/net13	vss	7.23918E-16
C1164	I0/I4049/net13	vss	7.44139E-16
C1165	I0/I2821/net13	vss	7.20083E-16
C1166	I0/I3302/net13	vss	7.20083E-16
C1167	I0/I3665/net13	vss	7.20083E-16
C1168	I0/I4059/net13	vss	7.42366E-16
C1169	I0/I5/net13	vss	7.23918E-16
C1170	I0/I3304/net13	vss	7.23918E-16
C1171	I0/I3675/net13	vss	7.23918E-16
C1172	I0/I4058/net13	vss	7.44139E-16
C1173	I0/I6/net13	vss	7.20083E-16
C1174	I0/I3289/net13	vss	7.20083E-16
C1175	I0/I3674/net13	vss	7.20083E-16
C1176	I0/I4066/net13	vss	7.42366E-16
C1177	I0/I82/net13	vss	7.23918E-16
C1178	I0/I3308/net13	vss	7.23918E-16
C1179	I0/I3682/net13	vss	7.23918E-16
C1180	I0/I4070/net13	vss	7.44139E-16
C1181	I0/I84/net13	vss	7.20313E-16
C1182	I0/I3283/net13	vss	7.20083E-16
C1183	I0/I3686/net13	vss	7.20083E-16
C1184	I0/I4072/net13	vss	7.42366E-16
C1185	I0/I3284/net13	vss	7.23918E-16
C1186	I0/I3688/net13	vss	7.23918E-16
C1187	I0/I4057/net13	vss	7.44139E-16
C1188	I0/I3292/net13	vss	7.20313E-16
C1189	I0/I3673/net13	vss	7.20083E-16
C1190	I0/I4076/net13	vss	7.42366E-16
C1191	I0/I3692/net13	vss	7.23918E-16
C1192	I0/I4051/net13	vss	7.44139E-16
C1193	I0/I3667/net13	vss	7.20083E-16
C1194	I0/I4052/net13	vss	7.42366E-16
C1195	I0/I3668/net13	vss	7.23918E-16
C1196	I0/I4060/net13	vss	7.35097E-16
C1197	I0/I3676/net13	vss	7.20313E-16
C1198	I33/net7	vss	1.15359E-15
C1199	I28/net7	vss	1.15048E-15
C1200	I0/I2807/net049	vss	9.09134E-16
C1201	I0/I2806/net049	vss	8.7256E-16
C1202	I0/I2817/net049	vss	8.95432E-16
C1203	I0/I2822/net049	vss	8.7256E-16
C1204	I0/I2818/net049	vss	8.95432E-16
C1205	I0/I3282/net049	vss	9.08793E-16
C1206	I0/I2814/net049	vss	8.7256E-16
C1207	I0/I3305/net049	vss	8.7222E-16
C1208	I0/I2815/net049	vss	8.95432E-16
C1209	I0/I3306/net049	vss	8.95091E-16
C1210	I0/I2819/net049	vss	8.7256E-16
C1211	I0/I4050/net049	vss	9.25916E-16
C1212	I0/I3295/net049	vss	8.7222E-16
C1213	I0/I2808/net049	vss	8.95432E-16
C1214	I0/I3666/net049	vss	9.08793E-16
C1215	I0/I4073/net049	vss	9.01201E-16
C1216	I0/I3309/net049	vss	8.95091E-16
C1217	I0/I2824/net049	vss	8.7256E-16
C1218	I0/I3689/net049	vss	8.7222E-16
C1219	I0/I4074/net049	vss	9.04706E-16
C1220	I0/I3297/net049	vss	8.7222E-16
C1221	I0/I2823/net049	vss	8.95432E-16
C1222	I0/I3690/net049	vss	8.95091E-16
C1223	I0/I4063/net049	vss	9.00873E-16
C1224	I0/I3293/net049	vss	8.95091E-16
C1225	I0/I2801/net049	vss	8.7256E-16
C1226	I0/I3679/net049	vss	8.7222E-16
C1227	I0/I4077/net049	vss	9.04706E-16
C1228	I0/I3299/net049	vss	8.7222E-16
C1229	I0/I2809/net049	vss	8.95432E-16
C1230	I0/I3693/net049	vss	8.95091E-16
C1231	I0/I4065/net049	vss	9.00873E-16
C1232	I0/I3285/net049	vss	8.95091E-16
C1233	I0/I2810/net049	vss	8.7256E-16
C1234	I0/I3681/net049	vss	8.7222E-16
C1235	I0/I4061/net049	vss	9.04706E-16
C1236	I0/I3296/net049	vss	8.7222E-16
C1237	I0/I2800/net049	vss	8.95432E-16
C1238	I0/I3677/net049	vss	8.95091E-16
C1239	I0/I4067/net049	vss	9.00873E-16
C1240	I0/I3294/net049	vss	8.95091E-16
C1241	I0/I2820/net049	vss	8.7256E-16
C1242	I0/I3683/net049	vss	8.7222E-16
C1243	I0/I4053/net049	vss	9.04706E-16
C1244	I0/I3288/net049	vss	8.7222E-16
C1245	I0/I2802/net049	vss	8.95432E-16
C1246	I0/I3669/net049	vss	8.95091E-16
C1247	I0/I4064/net049	vss	9.00873E-16
C1248	I0/I3286/net049	vss	8.95091E-16
C1249	I0/I2804/net049	vss	8.7256E-16
C1250	I0/I3279/net049	vss	8.7222E-16
C1251	I0/I3680/net049	vss	8.7222E-16
C1252	I0/I4062/net049	vss	9.04706E-16
C1253	I0/I2827/net049	vss	8.95432E-16
C1254	I0/I3278/net049	vss	8.95091E-16
C1255	I0/I3678/net049	vss	8.95091E-16
C1256	I0/I4056/net049	vss	9.00873E-16
C1257	I0/I2813/net049	vss	8.7256E-16
C1258	I0/I3300/net049	vss	8.7222E-16
C1259	I0/I3672/net049	vss	8.7222E-16
C1260	I0/I4054/net049	vss	9.04706E-16
C1261	I0/I2811/net049	vss	8.95432E-16
C1262	I0/I3303/net049	vss	8.95091E-16
C1263	I0/I3670/net049	vss	8.95091E-16
C1264	I0/I4047/net049	vss	9.00873E-16
C1265	I0/I2803/net049	vss	8.7256E-16
C1266	I0/I3280/net049	vss	8.7222E-16
C1267	I0/I3663/net049	vss	8.7222E-16
C1268	I0/I4046/net049	vss	9.04706E-16
C1269	I0/I2816/net049	vss	8.95432E-16
C1270	I0/I3287/net049	vss	8.95091E-16
C1271	I0/I3662/net049	vss	8.95091E-16
C1272	I0/I4068/net049	vss	9.00873E-16
C1273	I0/I2826/net049	vss	8.7256E-16
C1274	I0/I3301/net049	vss	8.7222E-16
C1275	I0/I3684/net049	vss	8.7222E-16
C1276	I0/I4071/net049	vss	9.04706E-16
C1277	I0/I2805/net049	vss	8.95432E-16
C1278	I0/I3307/net049	vss	8.95091E-16
C1279	I0/I3687/net049	vss	8.95091E-16
C1280	I0/I4048/net049	vss	9.00873E-16
C1281	I0/I2825/net049	vss	8.7256E-16
C1282	I0/I3281/net049	vss	8.7222E-16
C1283	I0/I3664/net049	vss	8.7222E-16
C1284	I0/I4055/net049	vss	9.04706E-16
C1285	I0/I2812/net049	vss	8.95432E-16
C1286	I0/I3291/net049	vss	8.95091E-16
C1287	I0/I3671/net049	vss	8.95091E-16
C1288	I0/I4069/net049	vss	9.00873E-16
C1289	I0/I2821/net049	vss	8.7256E-16
C1290	I0/I3290/net049	vss	8.7222E-16
C1291	I0/I3685/net049	vss	8.7222E-16
C1292	I0/I4075/net049	vss	9.04706E-16
C1293	I0/I5/net049	vss	8.95432E-16
C1294	I0/I3298/net049	vss	8.95091E-16
C1295	I0/I3691/net049	vss	8.95091E-16
C1296	I0/I4049/net049	vss	9.00873E-16
C1297	I0/I6/net049	vss	8.7256E-16
C1298	I0/I3302/net049	vss	8.7222E-16
C1299	I0/I3665/net049	vss	8.7222E-16
C1300	I0/I4059/net049	vss	9.04706E-16
C1301	I0/I82/net049	vss	8.95432E-16
C1302	I0/I3304/net049	vss	8.95091E-16
C1303	I0/I3675/net049	vss	8.95091E-16
C1304	I0/I4058/net049	vss	9.00873E-16
C1305	I0/I84/net049	vss	8.8E-16
C1306	I0/I3289/net049	vss	8.7222E-16
C1307	I0/I3674/net049	vss	8.7222E-16
C1308	I0/I4066/net049	vss	9.04706E-16
C1309	I0/I3308/net049	vss	8.95091E-16
C1310	I0/I3682/net049	vss	8.95091E-16
C1311	I0/I4070/net049	vss	9.00873E-16
C1312	I0/I3283/net049	vss	8.7222E-16
C1313	I0/I3686/net049	vss	8.7222E-16
C1314	I0/I4072/net049	vss	9.04706E-16
C1315	I0/I3284/net049	vss	8.95091E-16
C1316	I0/I3688/net049	vss	8.95091E-16
C1317	I0/I4057/net049	vss	9.00873E-16
C1318	I0/I3292/net049	vss	8.80256E-16
C1319	I0/I3673/net049	vss	8.7222E-16
C1320	I0/I4076/net049	vss	9.04706E-16
C1321	I0/I3692/net049	vss	8.95091E-16
C1322	I0/I4051/net049	vss	9.00873E-16
C1323	I0/I3667/net049	vss	8.7222E-16
C1324	I0/I4052/net049	vss	9.05034E-16
C1325	I3/net8	vss	7.85975E-16
C1326	I0/I3668/net049	vss	8.95091E-16
C1327	I0/I4060/net049	vss	8.98895E-16
C1328	I0/I3676/net049	vss	8.79659E-16
C1329	I33/net15	vss	1.16899E-15
C1330	I28/net15	vss	1.17914E-15
C1331	I0/I2863/net13	vss	7.29664E-16
C1332	I0/I2884/net13	vss	7.20083E-16
C1333	I0/I2878/net13	vss	7.23918E-16
C1334	I0/I2869/net13	vss	7.20083E-16
C1335	I0/I2870/net13	vss	7.23918E-16
C1336	I0/I2876/net13	vss	7.20083E-16
C1337	I0/I2873/net13	vss	7.23918E-16
C1338	I0/I3314/net13	vss	7.29664E-16
C1339	I0/I2882/net13	vss	7.20083E-16
C1340	I0/I4146/net13	vss	7.29091E-16
C1341	I0/I3337/net13	vss	7.20083E-16
C1342	I0/I2892/net13	vss	7.23918E-16
C1343	I0/I3698/net13	vss	7.29664E-16
C1344	I0/I4169/net13	vss	7.21505E-16
C1345	I0/I3338/net13	vss	7.23918E-16
C1346	I0/I2874/net13	vss	7.20083E-16
C1347	I0/I3721/net13	vss	7.20083E-16
C1348	I0/I4170/net13	vss	7.2534E-16
C1349	I0/I3327/net13	vss	7.20083E-16
C1350	I0/I2868/net13	vss	7.23918E-16
C1351	I0/I3722/net13	vss	7.23918E-16
C1352	I0/I4159/net13	vss	7.21505E-16
C1353	I0/I3341/net13	vss	7.23918E-16
C1354	I0/I2867/net13	vss	7.20083E-16
C1355	I0/I3711/net13	vss	7.20083E-16
C1356	I0/I4173/net13	vss	7.2534E-16
C1357	I0/I3329/net13	vss	7.20083E-16
C1358	I0/I2864/net13	vss	7.23918E-16
C1359	I0/I3725/net13	vss	7.23918E-16
C1360	I0/I4161/net13	vss	7.21505E-16
C1361	I0/I3325/net13	vss	7.23918E-16
C1362	I0/I2885/net13	vss	7.20083E-16
C1363	I0/I3713/net13	vss	7.20083E-16
C1364	I0/I4157/net13	vss	7.2534E-16
C1365	I0/I3331/net13	vss	7.20083E-16
C1366	I0/I2883/net13	vss	7.23918E-16
C1367	I0/I3709/net13	vss	7.23918E-16
C1368	I0/I4163/net13	vss	7.21505E-16
C1369	I0/I3317/net13	vss	7.23918E-16
C1370	I0/I2875/net13	vss	7.20083E-16
C1371	I0/I3715/net13	vss	7.20083E-16
C1372	I0/I4149/net13	vss	7.2534E-16
C1373	I0/I3328/net13	vss	7.20083E-16
C1374	I0/I2891/net13	vss	7.23918E-16
C1375	I0/I3701/net13	vss	7.23918E-16
C1376	I0/I4160/net13	vss	7.21505E-16
C1377	I0/I3326/net13	vss	7.23918E-16
C1378	I0/I2890/net13	vss	7.20083E-16
C1379	I0/I3712/net13	vss	7.20083E-16
C1380	I0/I4158/net13	vss	7.2534E-16
C1381	I0/I3320/net13	vss	7.20083E-16
C1382	I0/I2865/net13	vss	7.23918E-16
C1383	I0/I3710/net13	vss	7.23918E-16
C1384	I0/I4152/net13	vss	7.21505E-16
C1385	I0/I3318/net13	vss	7.23918E-16
C1386	I0/I2881/net13	vss	7.20083E-16
C1387	I0/I3704/net13	vss	7.20083E-16
C1388	I0/I4150/net13	vss	7.2534E-16
C1389	I0/I3311/net13	vss	7.20083E-16
C1390	I0/I2880/net13	vss	7.23918E-16
C1391	I0/I3702/net13	vss	7.23918E-16
C1392	I0/I4143/net13	vss	7.21505E-16
C1393	I0/I3310/net13	vss	7.23918E-16
C1394	I0/I2889/net13	vss	7.20083E-16
C1395	I0/I3695/net13	vss	7.20083E-16
C1396	I0/I4142/net13	vss	7.2534E-16
C1397	I0/I3332/net13	vss	7.20083E-16
C1398	I0/I2887/net13	vss	7.23918E-16
C1399	I0/I3694/net13	vss	7.23918E-16
C1400	I0/I4164/net13	vss	7.21505E-16
C1401	I0/I3335/net13	vss	7.23918E-16
C1402	I0/I2872/net13	vss	7.20083E-16
C1403	I0/I3716/net13	vss	7.20083E-16
C1404	I0/I4167/net13	vss	7.2534E-16
C1405	I0/I3312/net13	vss	7.20083E-16
C1406	I0/I2886/net13	vss	7.23918E-16
C1407	I0/I3719/net13	vss	7.23918E-16
C1408	I0/I4144/net13	vss	7.21505E-16
C1409	I0/I3319/net13	vss	7.23918E-16
C1410	I0/I2879/net13	vss	7.20083E-16
C1411	I0/I3696/net13	vss	7.20083E-16
C1412	I0/I4151/net13	vss	7.2534E-16
C1413	I0/I3333/net13	vss	7.20083E-16
C1414	I0/I2877/net13	vss	7.23918E-16
C1415	I0/I3703/net13	vss	7.23918E-16
C1416	I0/I4165/net13	vss	7.21505E-16
C1417	I0/I3339/net13	vss	7.23918E-16
C1418	I0/I2871/net13	vss	7.20083E-16
C1419	I0/I3717/net13	vss	7.20083E-16
C1420	I0/I4171/net13	vss	7.2534E-16
C1421	I0/I3313/net13	vss	7.20083E-16
C1422	I0/I2893/net13	vss	7.23918E-16
C1423	I0/I3723/net13	vss	7.23918E-16
C1424	I0/I4145/net13	vss	7.21505E-16
C1425	I0/I3323/net13	vss	7.23918E-16
C1426	I0/I2888/net13	vss	7.20083E-16
C1427	I0/I3697/net13	vss	7.20083E-16
C1428	I0/I4155/net13	vss	7.2534E-16
C1429	I0/I3322/net13	vss	7.20083E-16
C1430	I0/I2866/net13	vss	7.23918E-16
C1431	I0/I3707/net13	vss	7.23918E-16
C1432	I0/I4154/net13	vss	7.21505E-16
C1433	I0/I3330/net13	vss	7.23918E-16
C1434	I0/I2862/net13	vss	7.20313E-16
C1435	I0/I3706/net13	vss	7.20083E-16
C1436	I0/I4162/net13	vss	7.2534E-16
C1437	I0/I3334/net13	vss	7.20083E-16
C1438	I0/I3714/net13	vss	7.23918E-16
C1439	I0/I4166/net13	vss	7.21505E-16
C1440	I0/I3336/net13	vss	7.23918E-16
C1441	I0/I3718/net13	vss	7.20083E-16
C1442	I0/I4168/net13	vss	7.2534E-16
C1443	I0/I3321/net13	vss	7.20083E-16
C1444	I0/I3720/net13	vss	7.23918E-16
C1445	I0/I4153/net13	vss	7.21505E-16
C1446	I0/I3340/net13	vss	7.23918E-16
C1447	I0/I3705/net13	vss	7.20083E-16
C1448	I0/I4172/net13	vss	7.2534E-16
C1449	I0/I3315/net13	vss	7.20083E-16
C1450	I0/I3724/net13	vss	7.23918E-16
C1451	I0/I4147/net13	vss	7.21505E-16
C1452	I0/I3316/net13	vss	7.23918E-16
C1453	I0/I3699/net13	vss	7.20083E-16
C1454	I0/I4148/net13	vss	7.2534E-16
C1455	I0/I3324/net13	vss	7.20313E-16
C1456	I0/I3700/net13	vss	7.23918E-16
C1457	I0/I4156/net13	vss	7.19997E-16
C1458	I3/net20	vss	1.07252E-15
C1459	I0/I3708/net13	vss	7.20313E-16
C1460	I0/I2863/net049	vss	9.08034E-16
C1461	I0/I2884/net049	vss	8.71746E-16
C1462	I0/I2878/net049	vss	8.94618E-16
C1463	I0/I2869/net049	vss	8.71746E-16
C1464	I0/I2870/net049	vss	8.94618E-16
C1465	I0/I2876/net049	vss	8.71746E-16
C1466	I0/I2873/net049	vss	8.94618E-16
C1467	I0/I2882/net049	vss	8.71746E-16
C1468	I3/net23	vss	5.33607E-16
C1469	I0/I2892/net049	vss	8.94618E-16
C1470	I0/I3314/net049	vss	9.07863E-16
C1471	I0/I2874/net049	vss	8.71746E-16
C1472	I0/I4146/net049	vss	9.0756E-16
C1473	I0/I3337/net049	vss	8.71746E-16
C1474	I0/I2868/net049	vss	8.94618E-16
C1475	I0/I3698/net049	vss	9.08508E-16
C1476	I0/I4169/net049	vss	8.72084E-16
C1477	I0/I3338/net049	vss	8.94618E-16
C1478	I0/I2867/net049	vss	8.71746E-16
C1479	I0/I3721/net049	vss	8.7222E-16
C1480	I0/I4170/net049	vss	8.94956E-16
C1481	I0/I3327/net049	vss	8.71746E-16
C1482	I0/I2864/net049	vss	8.94618E-16
C1483	I0/I3722/net049	vss	8.95091E-16
C1484	I0/I4159/net049	vss	8.72084E-16
C1485	I0/I3341/net049	vss	8.94618E-16
C1486	I0/I2885/net049	vss	8.71746E-16
C1487	I0/I3711/net049	vss	8.7222E-16
C1488	I0/I4173/net049	vss	8.94956E-16
C1489	I0/I3329/net049	vss	8.71746E-16
C1490	I0/I2883/net049	vss	8.94618E-16
C1491	I0/I3725/net049	vss	8.95091E-16
C1492	I0/I4161/net049	vss	8.72084E-16
C1493	I0/I3325/net049	vss	8.94618E-16
C1494	I0/I2875/net049	vss	8.71746E-16
C1495	I0/I3713/net049	vss	8.7222E-16
C1496	I0/I4157/net049	vss	8.94956E-16
C1497	I0/I3331/net049	vss	8.71746E-16
C1498	I0/I2891/net049	vss	8.94618E-16
C1499	I0/I3709/net049	vss	8.95091E-16
C1500	I0/I4163/net049	vss	8.72084E-16
C1501	I0/I3317/net049	vss	8.94618E-16
C1502	I0/I2890/net049	vss	8.71746E-16
C1503	I0/I3715/net049	vss	8.7222E-16
C1504	I0/I4149/net049	vss	8.94956E-16
C1505	I0/I3328/net049	vss	8.71746E-16
C1506	I0/I2865/net049	vss	8.94618E-16
C1507	I0/I3701/net049	vss	8.95091E-16
C1508	I0/I4160/net049	vss	8.72084E-16
C1509	I0/I3326/net049	vss	8.94618E-16
C1510	I0/I2881/net049	vss	8.71746E-16
C1511	I0/I3712/net049	vss	8.7222E-16
C1512	I0/I4158/net049	vss	8.94956E-16
C1513	I0/I3320/net049	vss	8.71746E-16
C1514	I0/I2880/net049	vss	8.94618E-16
C1515	I0/I3710/net049	vss	8.95091E-16
C1516	I0/I4152/net049	vss	8.72084E-16
C1517	I0/I3318/net049	vss	8.94618E-16
C1518	I0/I2889/net049	vss	8.71746E-16
C1519	I0/I3704/net049	vss	8.7222E-16
C1520	I0/I4150/net049	vss	8.94956E-16
C1521	I0/I3311/net049	vss	8.71746E-16
C1522	I0/I2887/net049	vss	8.94618E-16
C1523	I0/I3702/net049	vss	8.95091E-16
C1524	I0/I4143/net049	vss	8.72084E-16
C1525	I0/I3310/net049	vss	8.94618E-16
C1526	I0/I2872/net049	vss	8.71746E-16
C1527	I0/I3695/net049	vss	8.7222E-16
C1528	I0/I4142/net049	vss	8.94956E-16
C1529	I0/I3332/net049	vss	8.71746E-16
C1530	I0/I2886/net049	vss	8.94618E-16
C1531	I0/I3694/net049	vss	8.95091E-16
C1532	I0/I4164/net049	vss	8.72084E-16
C1533	I0/I3335/net049	vss	8.94618E-16
C1534	I0/I2879/net049	vss	8.71746E-16
C1535	I0/I3716/net049	vss	8.7222E-16
C1536	I0/I4167/net049	vss	8.94956E-16
C1537	I0/I3312/net049	vss	8.71746E-16
C1538	I0/I2877/net049	vss	8.94618E-16
C1539	I0/I3719/net049	vss	8.95091E-16
C1540	I0/I4144/net049	vss	8.72084E-16
C1541	I0/I3319/net049	vss	8.94618E-16
C1542	I0/I2871/net049	vss	8.71746E-16
C1543	I0/I3696/net049	vss	8.7222E-16
C1544	I0/I4151/net049	vss	8.94956E-16
C1545	I0/I3333/net049	vss	8.71746E-16
C1546	I0/I2893/net049	vss	8.94618E-16
C1547	I0/I3703/net049	vss	8.95091E-16
C1548	I0/I4165/net049	vss	8.72084E-16
C1549	I0/I3339/net049	vss	8.94618E-16
C1550	I0/I2888/net049	vss	8.71746E-16
C1551	I0/I3717/net049	vss	8.7222E-16
C1552	I0/I4171/net049	vss	8.94956E-16
C1553	I0/I3313/net049	vss	8.71746E-16
C1554	I0/I2866/net049	vss	8.94618E-16
C1555	I0/I3723/net049	vss	8.95091E-16
C1556	I0/I4145/net049	vss	8.72084E-16
C1557	I0/I3323/net049	vss	8.94618E-16
C1558	I0/I2862/net049	vss	8.79783E-16
C1559	I0/I3697/net049	vss	8.7222E-16
C1560	I0/I4155/net049	vss	8.94956E-16
C1561	I0/I3322/net049	vss	8.71746E-16
C1562	I0/I3707/net049	vss	8.95091E-16
C1563	I0/I4154/net049	vss	8.72084E-16
C1564	I0/I3330/net049	vss	8.94618E-16
C1565	I0/I3706/net049	vss	8.7222E-16
C1566	I0/I4162/net049	vss	8.94956E-16
C1567	I0/I3334/net049	vss	8.71746E-16
C1568	I0/I3714/net049	vss	8.95091E-16
C1569	I0/I4166/net049	vss	8.72084E-16
C1570	I0/I3336/net049	vss	8.94618E-16
C1571	I0/I3718/net049	vss	8.7222E-16
C1572	I0/I4168/net049	vss	8.94956E-16
C1573	I0/I3321/net049	vss	8.71746E-16
C1574	I0/I3720/net049	vss	8.95091E-16
C1575	I0/I4153/net049	vss	8.72084E-16
C1576	I0/I3340/net049	vss	8.94618E-16
C1577	I0/I3705/net049	vss	8.7222E-16
C1578	I0/I4172/net049	vss	8.94956E-16
C1579	I0/I3315/net049	vss	8.71746E-16
C1580	I0/I3724/net049	vss	8.95091E-16
C1581	I0/I4147/net049	vss	8.72084E-16
C1582	I0/I3316/net049	vss	8.94618E-16
C1583	I0/I3699/net049	vss	8.7222E-16
C1584	I0/I4148/net049	vss	8.94956E-16
C1585	I0/I3324/net049	vss	8.79783E-16
C1586	I0/I3700/net049	vss	8.95091E-16
C1587	I0/I4156/net049	vss	8.79526E-16
C1588	I3/net24	vss	6.07779E-16
C1589	I0/I3708/net049	vss	8.79659E-16
C1590	I116/net0113	vss	3.31689E-15
C1591	I11/net8	vss	8.24248E-16
C1592	I6/net8	vss	7.88173E-16
C1593	I0/I2925/net13	vss	7.29837E-16
C1594	I0/I2904/net13	vss	7.20083E-16
C1595	I0/I2900/net13	vss	7.23918E-16
C1596	I0/I2899/net13	vss	7.20083E-16
C1597	I0/I2898/net13	vss	7.23918E-16
C1598	I0/I2911/net13	vss	7.20083E-16
C1599	I0/I3346/net13	vss	7.29699E-16
C1600	I0/I2921/net13	vss	7.23918E-16
C1601	I0/I3369/net13	vss	7.20083E-16
C1602	I0/I2924/net13	vss	7.20083E-16
C1603	I0/I3370/net13	vss	7.23918E-16
C1604	I0/I2917/net13	vss	7.23918E-16
C1605	I0/I4178/net13	vss	7.29983E-16
C1606	I0/I3359/net13	vss	7.20083E-16
C1607	I0/I2907/net13	vss	7.20083E-16
C1608	I0/I4201/net13	vss	7.20083E-16
C1609	I0/I3373/net13	vss	7.23918E-16
C1610	I0/I2897/net13	vss	7.23918E-16
C1611	I0/I3730/net13	vss	7.29837E-16
C1612	I0/I4202/net13	vss	7.23918E-16
C1613	I0/I3361/net13	vss	7.20083E-16
C1614	I0/I2896/net13	vss	7.20083E-16
C1615	I0/I3753/net13	vss	7.20083E-16
C1616	I0/I4191/net13	vss	7.20083E-16
C1617	I0/I3357/net13	vss	7.23918E-16
C1618	I0/I2916/net13	vss	7.23918E-16
C1619	I0/I3754/net13	vss	7.23918E-16
C1620	I0/I4205/net13	vss	7.23918E-16
C1621	I0/I3363/net13	vss	7.20083E-16
C1622	I0/I2906/net13	vss	7.20083E-16
C1623	I0/I3743/net13	vss	7.20083E-16
C1624	I0/I4193/net13	vss	7.20083E-16
C1625	I0/I3349/net13	vss	7.23918E-16
C1626	I0/I2918/net13	vss	7.23918E-16
C1627	I0/I3757/net13	vss	7.23918E-16
C1628	I0/I4189/net13	vss	7.23918E-16
C1629	I0/I3360/net13	vss	7.20083E-16
C1630	I0/I2912/net13	vss	7.20083E-16
C1631	I0/I3745/net13	vss	7.20083E-16
C1632	I0/I4195/net13	vss	7.20083E-16
C1633	I0/I3358/net13	vss	7.23918E-16
C1634	I0/I2908/net13	vss	7.23918E-16
C1635	I0/I3741/net13	vss	7.23918E-16
C1636	I0/I4181/net13	vss	7.23918E-16
C1637	I0/I3352/net13	vss	7.20083E-16
C1638	I0/I2913/net13	vss	7.20083E-16
C1639	I0/I3747/net13	vss	7.20083E-16
C1640	I0/I4192/net13	vss	7.20083E-16
C1641	I0/I3350/net13	vss	7.23918E-16
C1642	I0/I2914/net13	vss	7.23918E-16
C1643	I0/I3733/net13	vss	7.23918E-16
C1644	I0/I4190/net13	vss	7.23918E-16
C1645	I0/I3343/net13	vss	7.20083E-16
C1646	I0/I2901/net13	vss	7.20083E-16
C1647	I0/I3744/net13	vss	7.20083E-16
C1648	I0/I4184/net13	vss	7.20083E-16
C1649	I0/I3342/net13	vss	7.23918E-16
C1650	I0/I2902/net13	vss	7.23918E-16
C1651	I0/I3742/net13	vss	7.23918E-16
C1652	I0/I4182/net13	vss	7.23918E-16
C1653	I0/I3364/net13	vss	7.20083E-16
C1654	I0/I2915/net13	vss	7.20083E-16
C1655	I0/I3736/net13	vss	7.20083E-16
C1656	I0/I4175/net13	vss	7.20083E-16
C1657	I0/I3367/net13	vss	7.23918E-16
C1658	I0/I2920/net13	vss	7.23918E-16
C1659	I0/I3734/net13	vss	7.23918E-16
C1660	I0/I4174/net13	vss	7.23918E-16
C1661	I0/I3344/net13	vss	7.20083E-16
C1662	I0/I2905/net13	vss	7.20083E-16
C1663	I0/I3727/net13	vss	7.20083E-16
C1664	I0/I4196/net13	vss	7.20083E-16
C1665	I0/I3351/net13	vss	7.23918E-16
C1666	I0/I2910/net13	vss	7.23918E-16
C1667	I0/I3726/net13	vss	7.23918E-16
C1668	I0/I4199/net13	vss	7.23918E-16
C1669	I0/I3365/net13	vss	7.20083E-16
C1670	I0/I2919/net13	vss	7.20083E-16
C1671	I0/I3748/net13	vss	7.20083E-16
C1672	I0/I4176/net13	vss	7.20083E-16
C1673	I0/I3371/net13	vss	7.23918E-16
C1674	I0/I2922/net13	vss	7.23918E-16
C1675	I0/I3751/net13	vss	7.23918E-16
C1676	I0/I4183/net13	vss	7.23918E-16
C1677	I0/I3345/net13	vss	7.20083E-16
C1678	I0/I2903/net13	vss	7.20083E-16
C1679	I0/I3728/net13	vss	7.20083E-16
C1680	I0/I4197/net13	vss	7.20083E-16
C1681	I0/I3355/net13	vss	7.23918E-16
C1682	I0/I2923/net13	vss	7.23918E-16
C1683	I0/I3735/net13	vss	7.23918E-16
C1684	I0/I4203/net13	vss	7.23918E-16
C1685	I0/I3354/net13	vss	7.20083E-16
C1686	I0/I2909/net13	vss	7.20083E-16
C1687	I0/I3749/net13	vss	7.20083E-16
C1688	I0/I4177/net13	vss	7.20083E-16
C1689	I0/I3362/net13	vss	7.23918E-16
C1690	I0/I2895/net13	vss	7.23918E-16
C1691	I0/I3755/net13	vss	7.23918E-16
C1692	I0/I4187/net13	vss	7.23918E-16
C1693	I0/I3366/net13	vss	7.20083E-16
C1694	I0/I2894/net13	vss	7.20313E-16
C1695	I0/I3729/net13	vss	7.20083E-16
C1696	I0/I4186/net13	vss	7.20083E-16
C1697	I0/I3368/net13	vss	7.23918E-16
C1698	I0/I3739/net13	vss	7.23918E-16
C1699	I0/I4194/net13	vss	7.23918E-16
C1700	I0/I3353/net13	vss	7.20083E-16
C1701	I0/I3738/net13	vss	7.20083E-16
C1702	I0/I4198/net13	vss	7.20083E-16
C1703	I0/I3372/net13	vss	7.23918E-16
C1704	I0/I3746/net13	vss	7.23918E-16
C1705	I0/I4200/net13	vss	7.23918E-16
C1706	I0/I3347/net13	vss	7.20083E-16
C1707	I0/I3750/net13	vss	7.20083E-16
C1708	I0/I4185/net13	vss	7.20083E-16
C1709	I0/I3348/net13	vss	7.23918E-16
C1710	I0/I3752/net13	vss	7.23918E-16
C1711	I0/I4204/net13	vss	7.23918E-16
C1712	I0/I3356/net13	vss	7.20313E-16
C1713	I0/I3737/net13	vss	7.20083E-16
C1714	I0/I4179/net13	vss	7.20083E-16
C1715	I0/I3756/net13	vss	7.23918E-16
C1716	I0/I4180/net13	vss	7.23918E-16
C1717	I0/I3731/net13	vss	7.20083E-16
C1718	I0/I4188/net13	vss	7.20313E-16
C1719	I0/I3732/net13	vss	7.23918E-16
C1720	I0/I3740/net13	vss	7.20313E-16
C1721	I0/I2925/net049	vss	9.09689E-16
C1722	I0/I2904/net049	vss	8.71746E-16
C1723	I0/I2900/net049	vss	8.94618E-16
C1724	I0/I2899/net049	vss	8.71746E-16
C1725	I0/I2898/net049	vss	8.94618E-16
C1726	I0/I2911/net049	vss	8.71746E-16
C1727	I0/I2921/net049	vss	8.94618E-16
C1728	I24/net7	vss	1.16419E-15
C1729	I0/I2924/net049	vss	8.71746E-16
C1730	I0/I2917/net049	vss	8.94618E-16
C1731	I0/I2907/net049	vss	8.71746E-16
C1732	I11/net20	vss	1.07324E-15
C1733	I0/I3346/net049	vss	9.09518E-16
C1734	I0/I2897/net049	vss	8.94618E-16
C1735	I6/net20	vss	1.07039E-15
C1736	I0/I4178/net049	vss	9.09801E-16
C1737	I0/I3369/net049	vss	8.71746E-16
C1738	I0/I2896/net049	vss	8.71746E-16
C1739	I6/net23	vss	5.3506E-16
C1740	I0/I4201/net049	vss	8.71746E-16
C1741	I0/I3370/net049	vss	8.94618E-16
C1742	I0/I2916/net049	vss	8.94618E-16
C1743	I0/I3730/net049	vss	9.09689E-16
C1744	I0/I4202/net049	vss	8.94618E-16
C1745	I0/I3359/net049	vss	8.71746E-16
C1746	I0/I2906/net049	vss	8.71746E-16
C1747	I0/I3753/net049	vss	8.71746E-16
C1748	I0/I4191/net049	vss	8.71746E-16
C1749	I0/I3373/net049	vss	8.94618E-16
C1750	I0/I2918/net049	vss	8.94618E-16
C1751	I0/I3754/net049	vss	8.94618E-16
C1752	I0/I4205/net049	vss	8.94618E-16
C1753	I0/I3361/net049	vss	8.71746E-16
C1754	I0/I2912/net049	vss	8.71746E-16
C1755	I0/I3743/net049	vss	8.71746E-16
C1756	I0/I4193/net049	vss	8.71746E-16
C1757	I0/I3357/net049	vss	8.94618E-16
C1758	I0/I2908/net049	vss	8.94618E-16
C1759	I0/I3757/net049	vss	8.94618E-16
C1760	I0/I4189/net049	vss	8.94618E-16
C1761	I0/I3363/net049	vss	8.71746E-16
C1762	I0/I2913/net049	vss	8.71746E-16
C1763	I0/I3745/net049	vss	8.71746E-16
C1764	I0/I4195/net049	vss	8.71746E-16
C1765	I0/I3349/net049	vss	8.94618E-16
C1766	I0/I2914/net049	vss	8.94618E-16
C1767	I0/I3741/net049	vss	8.94618E-16
C1768	I0/I4181/net049	vss	8.94618E-16
C1769	I0/I3360/net049	vss	8.71746E-16
C1770	I0/I2901/net049	vss	8.71746E-16
C1771	I0/I3747/net049	vss	8.71746E-16
C1772	I0/I4192/net049	vss	8.71746E-16
C1773	I0/I3358/net049	vss	8.94618E-16
C1774	I0/I2902/net049	vss	8.94618E-16
C1775	I0/I3733/net049	vss	8.94618E-16
C1776	I0/I4190/net049	vss	8.94618E-16
C1777	I0/I3352/net049	vss	8.71746E-16
C1778	I0/I2915/net049	vss	8.71746E-16
C1779	I0/I3744/net049	vss	8.71746E-16
C1780	I0/I4184/net049	vss	8.71746E-16
C1781	I0/I3350/net049	vss	8.94618E-16
C1782	I0/I2920/net049	vss	8.94618E-16
C1783	I0/I3742/net049	vss	8.94618E-16
C1784	I0/I4182/net049	vss	8.94618E-16
C1785	I0/I3343/net049	vss	8.71746E-16
C1786	I0/I2905/net049	vss	8.71746E-16
C1787	I0/I3736/net049	vss	8.71746E-16
C1788	I0/I4175/net049	vss	8.71746E-16
C1789	I0/I3342/net049	vss	8.94618E-16
C1790	I0/I2910/net049	vss	8.94618E-16
C1791	I0/I3734/net049	vss	8.94618E-16
C1792	I0/I4174/net049	vss	8.94618E-16
C1793	I0/I3364/net049	vss	8.71746E-16
C1794	I0/I2919/net049	vss	8.71746E-16
C1795	I0/I3727/net049	vss	8.71746E-16
C1796	I0/I4196/net049	vss	8.71746E-16
C1797	I0/I3367/net049	vss	8.94618E-16
C1798	I0/I2922/net049	vss	8.94618E-16
C1799	I0/I3726/net049	vss	8.94618E-16
C1800	I0/I4199/net049	vss	8.94618E-16
C1801	I0/I3344/net049	vss	8.71746E-16
C1802	I0/I2903/net049	vss	8.71746E-16
C1803	I0/I3748/net049	vss	8.71746E-16
C1804	I0/I4176/net049	vss	8.71746E-16
C1805	I0/I3351/net049	vss	8.94618E-16
C1806	I0/I2923/net049	vss	8.94618E-16
C1807	I0/I3751/net049	vss	8.94618E-16
C1808	I0/I4183/net049	vss	8.94618E-16
C1809	I0/I3365/net049	vss	8.71746E-16
C1810	I0/I2909/net049	vss	8.71746E-16
C1811	I0/I3728/net049	vss	8.71746E-16
C1812	I0/I4197/net049	vss	8.71746E-16
C1813	I0/I3371/net049	vss	8.94618E-16
C1814	I0/I2895/net049	vss	8.94618E-16
C1815	I0/I3735/net049	vss	8.94618E-16
C1816	I0/I4203/net049	vss	8.94618E-16
C1817	I0/I3345/net049	vss	8.71746E-16
C1818	I0/I2894/net049	vss	8.79186E-16
C1819	I0/I3749/net049	vss	8.71746E-16
C1820	I0/I4177/net049	vss	8.71746E-16
C1821	I0/I3355/net049	vss	8.94618E-16
C1822	I0/I3755/net049	vss	8.94618E-16
C1823	I0/I4187/net049	vss	8.94618E-16
C1824	I0/I3354/net049	vss	8.71746E-16
C1825	I116/net0125	vss	3.32453E-15
C1826	I0/I3729/net049	vss	8.71746E-16
C1827	I0/I4186/net049	vss	8.71746E-16
C1828	I0/I3362/net049	vss	8.94618E-16
C1829	I0/I3739/net049	vss	8.94618E-16
C1830	I0/I4194/net049	vss	8.94618E-16
C1831	I0/I3366/net049	vss	8.71746E-16
C1832	I0/I3738/net049	vss	8.71746E-16
C1833	I0/I4198/net049	vss	8.71746E-16
C1834	I0/I3368/net049	vss	8.94618E-16
C1835	I0/I3746/net049	vss	8.94618E-16
C1836	I0/I4200/net049	vss	8.94618E-16
C1837	I0/I3353/net049	vss	8.71746E-16
C1838	I0/I3750/net049	vss	8.71746E-16
C1839	I0/I4185/net049	vss	8.71746E-16
C1840	I0/I3372/net049	vss	8.94618E-16
C1841	I0/I3752/net049	vss	8.94618E-16
C1842	I0/I4204/net049	vss	8.94618E-16
C1843	I0/I3347/net049	vss	8.71746E-16
C1844	I0/I3737/net049	vss	8.71746E-16
C1845	I0/I4179/net049	vss	8.71746E-16
C1846	I0/I3348/net049	vss	8.94618E-16
C1847	I0/I3756/net049	vss	8.94618E-16
C1848	I0/I4180/net049	vss	8.94618E-16
C1849	I0/I3356/net049	vss	8.79186E-16
C1850	I0/I3731/net049	vss	8.71746E-16
C1851	I0/I4188/net049	vss	8.79783E-16
C1852	I0/I3732/net049	vss	8.94618E-16
C1853	I0/I3740/net049	vss	8.79186E-16
C1854	I11/net23	vss	5.29607E-16
C1855	I6/net24	vss	6.80415E-16
C1856	I24/net15	vss	1.17186E-15
C1857	I11/net24	vss	7.14538E-16
C1858	I0/I2937/net13	vss	7.34169E-16
C1859	I0/I2939/net13	vss	7.24349E-16
C1860	I0/I2927/net13	vss	7.27551E-16
C1861	I0/I2931/net13	vss	7.23621E-16
C1862	I0/I2930/net13	vss	7.27699E-16
C1863	I0/I2944/net13	vss	7.23406E-16
C1864	I0/I2946/net13	vss	7.27466E-16
C1865	I0/I2955/net13	vss	7.22013E-16
C1866	I0/I2954/net13	vss	7.27272E-16
C1867	I0/I2945/net13	vss	7.22078E-16
C1868	I0/I2929/net13	vss	7.2733E-16
C1869	I0/I2928/net13	vss	7.21695E-16
C1870	I0/I4210/net13	vss	7.30111E-16
C1871	I0/I2932/net13	vss	7.27192E-16
C1872	I0/I3762/net13	vss	7.29973E-16
C1873	I0/I4233/net13	vss	7.20083E-16
C1874	I0/I3378/net13	vss	7.29973E-16
C1875	I0/I2942/net13	vss	7.22024E-16
C1876	I0/I3785/net13	vss	7.20083E-16
C1877	I0/I4234/net13	vss	7.23918E-16
C1878	I0/I3401/net13	vss	7.20083E-16
C1879	I0/I2952/net13	vss	7.27094E-16
C1880	I0/I3786/net13	vss	7.23918E-16
C1881	I0/I4223/net13	vss	7.20083E-16
C1882	I0/I3402/net13	vss	7.23918E-16
C1883	I0/I2948/net13	vss	7.21709E-16
C1884	I0/I3775/net13	vss	7.20083E-16
C1885	I0/I4237/net13	vss	7.23918E-16
C1886	I0/I3391/net13	vss	7.20083E-16
C1887	I0/I2943/net13	vss	7.24787E-16
C1888	I0/I3789/net13	vss	7.23918E-16
C1889	I0/I4225/net13	vss	7.20083E-16
C1890	I0/I3405/net13	vss	7.23918E-16
C1891	I0/I2950/net13	vss	7.21648E-16
C1892	I0/I3777/net13	vss	7.20083E-16
C1893	I0/I4221/net13	vss	7.23918E-16
C1894	I0/I3393/net13	vss	7.20083E-16
C1895	I0/I2947/net13	vss	7.24511E-16
C1896	I0/I3773/net13	vss	7.23918E-16
C1897	I0/I4227/net13	vss	7.20083E-16
C1898	I0/I3389/net13	vss	7.23918E-16
C1899	I0/I2935/net13	vss	7.21722E-16
C1900	I0/I3779/net13	vss	7.20083E-16
C1901	I0/I4213/net13	vss	7.23918E-16
C1902	I0/I3395/net13	vss	7.20083E-16
C1903	I0/I2938/net13	vss	7.24666E-16
C1904	I0/I3765/net13	vss	7.23918E-16
C1905	I0/I4224/net13	vss	7.20083E-16
C1906	I0/I3381/net13	vss	7.23918E-16
C1907	I0/I2949/net13	vss	7.21694E-16
C1908	I0/I3776/net13	vss	7.20083E-16
C1909	I0/I4222/net13	vss	7.23918E-16
C1910	I0/I3392/net13	vss	7.20083E-16
C1911	I0/I2953/net13	vss	7.2449E-16
C1912	I0/I3774/net13	vss	7.23918E-16
C1913	I0/I4216/net13	vss	7.20083E-16
C1914	I0/I3390/net13	vss	7.23918E-16
C1915	I0/I2941/net13	vss	7.21901E-16
C1916	I0/I3768/net13	vss	7.20083E-16
C1917	I0/I4214/net13	vss	7.23918E-16
C1918	I0/I3384/net13	vss	7.20083E-16
C1919	I0/I2936/net13	vss	7.24944E-16
C1920	I0/I3766/net13	vss	7.23918E-16
C1921	I0/I4207/net13	vss	7.20083E-16
C1922	I0/I3382/net13	vss	7.23918E-16
C1923	I0/I2957/net13	vss	7.21851E-16
C1924	I0/I3759/net13	vss	7.20083E-16
C1925	I0/I4206/net13	vss	7.23918E-16
C1926	I0/I3375/net13	vss	7.20083E-16
C1927	I0/I2956/net13	vss	7.24797E-16
C1928	I0/I3758/net13	vss	7.23918E-16
C1929	I0/I4228/net13	vss	7.20083E-16
C1930	I0/I3374/net13	vss	7.23918E-16
C1931	I0/I2940/net13	vss	7.21879E-16
C1932	I0/I3780/net13	vss	7.20083E-16
C1933	I0/I4231/net13	vss	7.23918E-16
C1934	I0/I3396/net13	vss	7.20083E-16
C1935	I0/I2951/net13	vss	7.25498E-16
C1936	I0/I3783/net13	vss	7.23918E-16
C1937	I0/I4208/net13	vss	7.20083E-16
C1938	I0/I3399/net13	vss	7.23918E-16
C1939	I0/I2933/net13	vss	7.22101E-16
C1940	I0/I3760/net13	vss	7.20083E-16
C1941	I0/I4215/net13	vss	7.23918E-16
C1942	I0/I3376/net13	vss	7.20083E-16
C1943	I0/I2934/net13	vss	7.24849E-16
C1944	I0/I3767/net13	vss	7.23918E-16
C1945	I0/I4229/net13	vss	7.20083E-16
C1946	I0/I3383/net13	vss	7.23918E-16
C1947	I0/I2926/net13	vss	7.21836E-16
C1948	I0/I3781/net13	vss	7.20083E-16
C1949	I0/I4235/net13	vss	7.23918E-16
C1950	I0/I3397/net13	vss	7.20083E-16
C1951	I0/I3787/net13	vss	7.23918E-16
C1952	I0/I4209/net13	vss	7.20083E-16
C1953	I0/I3403/net13	vss	7.23918E-16
C1954	I0/I3761/net13	vss	7.20083E-16
C1955	I0/I4219/net13	vss	7.23918E-16
C1956	I0/I3377/net13	vss	7.20083E-16
C1957	I0/I3771/net13	vss	7.23918E-16
C1958	I0/I4218/net13	vss	7.20083E-16
C1959	I0/I3387/net13	vss	7.23918E-16
C1960	I0/I3770/net13	vss	7.20083E-16
C1961	I0/I4226/net13	vss	7.23918E-16
C1962	I0/I3386/net13	vss	7.20083E-16
C1963	I0/I3778/net13	vss	7.23918E-16
C1964	I0/I4230/net13	vss	7.20083E-16
C1965	I0/I3394/net13	vss	7.23918E-16
C1966	I0/I3782/net13	vss	7.20083E-16
C1967	I0/I4232/net13	vss	7.23918E-16
C1968	I0/I3398/net13	vss	7.20083E-16
C1969	I0/I3784/net13	vss	7.23918E-16
C1970	I0/I4217/net13	vss	7.20083E-16
C1971	I0/I3400/net13	vss	7.23918E-16
C1972	I0/I3769/net13	vss	7.20083E-16
C1973	I0/I4236/net13	vss	7.23918E-16
C1974	I0/I3385/net13	vss	7.20083E-16
C1975	I0/I3788/net13	vss	7.23918E-16
C1976	I0/I4211/net13	vss	7.20083E-16
C1977	I0/I3404/net13	vss	7.23918E-16
C1978	I0/I3763/net13	vss	7.20083E-16
C1979	I0/I4212/net13	vss	7.23918E-16
C1980	I0/I3379/net13	vss	7.20083E-16
C1981	I0/I3764/net13	vss	7.23918E-16
C1982	I0/I4220/net13	vss	7.20313E-16
C1983	I0/I3380/net13	vss	7.23918E-16
C1984	I0/I3772/net13	vss	7.20313E-16
C1985	I32/net7	vss	1.152E-15
C1986	I0/I3388/net13	vss	7.20313E-16
C1987	I27/net7	vss	1.15232E-15
C1988	I0/I2937/net049	vss	9.04908E-16
C1989	I0/I2939/net049	vss	8.68918E-16
C1990	I0/I2927/net049	vss	8.90834E-16
C1991	I0/I2931/net049	vss	8.71198E-16
C1992	I0/I2930/net049	vss	8.9021E-16
C1993	I0/I2944/net049	vss	8.64443E-16
C1994	I0/I2946/net049	vss	8.90155E-16
C1995	I0/I2955/net049	vss	8.67955E-16
C1996	I0/I2954/net049	vss	8.89832E-16
C1997	I0/I2945/net049	vss	8.67592E-16
C1998	I0/I2929/net049	vss	8.90866E-16
C1999	I0/I2928/net049	vss	8.66948E-16
C2000	I0/I2932/net049	vss	8.92019E-16
C2001	I0/I2942/net049	vss	8.68667E-16
C2002	I0/I4210/net049	vss	9.08532E-16
C2003	I0/I2952/net049	vss	8.88956E-16
C2004	I0/I3762/net049	vss	9.08701E-16
C2005	I0/I4233/net049	vss	8.7222E-16
C2006	I0/I3378/net049	vss	9.07887E-16
C2007	I0/I2948/net049	vss	8.73525E-16
C2008	I0/I3785/net049	vss	8.7256E-16
C2009	I0/I4234/net049	vss	8.95091E-16
C2010	I0/I3401/net049	vss	8.71746E-16
C2011	I0/I2943/net049	vss	8.94111E-16
C2012	I0/I3786/net049	vss	8.95432E-16
C2013	I0/I4223/net049	vss	8.7222E-16
C2014	I0/I3402/net049	vss	8.94618E-16
C2015	I0/I2950/net049	vss	8.70584E-16
C2016	I0/I3775/net049	vss	8.7256E-16
C2017	I0/I4237/net049	vss	8.95091E-16
C2018	I0/I3391/net049	vss	8.71746E-16
C2019	I0/I2947/net049	vss	8.94409E-16
C2020	I0/I3789/net049	vss	8.95432E-16
C2021	I0/I4225/net049	vss	8.7222E-16
C2022	I0/I3405/net049	vss	8.94618E-16
C2023	I0/I2935/net049	vss	8.67507E-16
C2024	I0/I3777/net049	vss	8.7256E-16
C2025	I0/I4221/net049	vss	8.95091E-16
C2026	I0/I3393/net049	vss	8.71746E-16
C2027	I0/I2938/net049	vss	8.90145E-16
C2028	I0/I3773/net049	vss	8.95432E-16
C2029	I0/I4227/net049	vss	8.7222E-16
C2030	I0/I3389/net049	vss	8.94618E-16
C2031	I0/I2949/net049	vss	8.6975E-16
C2032	I0/I3779/net049	vss	8.7256E-16
C2033	I0/I4213/net049	vss	8.95091E-16
C2034	I0/I3395/net049	vss	8.71746E-16
C2035	I0/I2953/net049	vss	8.90205E-16
C2036	I0/I3765/net049	vss	8.95432E-16
C2037	I0/I4224/net049	vss	8.7222E-16
C2038	I0/I3381/net049	vss	8.94618E-16
C2039	I0/I2941/net049	vss	8.6873E-16
C2040	I0/I3776/net049	vss	8.7256E-16
C2041	I0/I4222/net049	vss	8.95091E-16
C2042	I0/I3392/net049	vss	8.71746E-16
C2043	I0/I2936/net049	vss	8.89869E-16
C2044	I0/I3774/net049	vss	8.95432E-16
C2045	I0/I4216/net049	vss	8.7222E-16
C2046	I0/I3390/net049	vss	8.94618E-16
C2047	I0/I2957/net049	vss	8.69528E-16
C2048	I0/I3768/net049	vss	8.7256E-16
C2049	I0/I4214/net049	vss	8.95091E-16
C2050	I0/I3384/net049	vss	8.71746E-16
C2051	I0/I2956/net049	vss	8.89941E-16
C2052	I0/I3766/net049	vss	8.95432E-16
C2053	I0/I4207/net049	vss	8.7222E-16
C2054	I0/I3382/net049	vss	8.94618E-16
C2055	I0/I2940/net049	vss	8.72669E-16
C2056	I0/I3759/net049	vss	8.7256E-16
C2057	I0/I4206/net049	vss	8.95091E-16
C2058	I0/I3375/net049	vss	8.71746E-16
C2059	I0/I2951/net049	vss	8.91705E-16
C2060	I0/I3758/net049	vss	8.95432E-16
C2061	I0/I4228/net049	vss	8.7222E-16
C2062	I0/I3374/net049	vss	8.94618E-16
C2063	I0/I2933/net049	vss	8.6437E-16
C2064	I0/I3780/net049	vss	8.7256E-16
C2065	I0/I4231/net049	vss	8.95091E-16
C2066	I0/I3396/net049	vss	8.71746E-16
C2067	I0/I2934/net049	vss	8.90674E-16
C2068	I0/I3783/net049	vss	8.95432E-16
C2069	I0/I4208/net049	vss	8.7222E-16
C2070	I0/I3399/net049	vss	8.94618E-16
C2071	I0/I2926/net049	vss	8.75844E-16
C2072	I0/I3760/net049	vss	8.7256E-16
C2073	I0/I4215/net049	vss	8.95091E-16
C2074	I0/I3376/net049	vss	8.71746E-16
C2075	I0/I3767/net049	vss	8.95432E-16
C2076	I0/I4229/net049	vss	8.7222E-16
C2077	I0/I3383/net049	vss	8.94618E-16
C2078	I0/I3781/net049	vss	8.7256E-16
C2079	I0/I4235/net049	vss	8.95091E-16
C2080	I0/I3397/net049	vss	8.71746E-16
C2081	I0/I3787/net049	vss	8.95432E-16
C2082	I0/I4209/net049	vss	8.7222E-16
C2083	I0/I3403/net049	vss	8.94618E-16
C2084	I0/I3761/net049	vss	8.7256E-16
C2085	I0/I4219/net049	vss	8.95091E-16
C2086	I0/I3377/net049	vss	8.71746E-16
C2087	I0/I3771/net049	vss	8.95432E-16
C2088	I0/I4218/net049	vss	8.7222E-16
C2089	I0/I3387/net049	vss	8.94618E-16
C2090	I0/I3770/net049	vss	8.7256E-16
C2091	I0/I4226/net049	vss	8.95091E-16
C2092	I0/I3386/net049	vss	8.71746E-16
C2093	I0/I3778/net049	vss	8.95432E-16
C2094	I0/I4230/net049	vss	8.7222E-16
C2095	I0/I3394/net049	vss	8.94618E-16
C2096	I0/I3782/net049	vss	8.7256E-16
C2097	I0/I4232/net049	vss	8.95091E-16
C2098	I0/I3398/net049	vss	8.71746E-16
C2099	I0/I3784/net049	vss	8.95432E-16
C2100	I0/I4217/net049	vss	8.7222E-16
C2101	I0/I3400/net049	vss	8.94618E-16
C2102	I0/I3769/net049	vss	8.7256E-16
C2103	I0/I4236/net049	vss	8.95091E-16
C2104	I0/I3385/net049	vss	8.71746E-16
C2105	I0/I3788/net049	vss	8.95432E-16
C2106	I0/I4211/net049	vss	8.7222E-16
C2107	I0/I3404/net049	vss	8.94618E-16
C2108	I0/I3763/net049	vss	8.7256E-16
C2109	I0/I4212/net049	vss	8.95091E-16
C2110	I0/I3379/net049	vss	8.71746E-16
C2111	I0/I3764/net049	vss	8.95432E-16
C2112	I0/I4220/net049	vss	8.79659E-16
C2113	I0/I3380/net049	vss	8.94618E-16
C2114	I0/I3772/net049	vss	8.8E-16
C2115	I0/I3388/net049	vss	8.79783E-16
C2116	I27/net15	vss	1.18047E-15
C2117	I32/net15	vss	1.18544E-15
C2118	I116/net0133	vss	2.18651E-15
C2119	I2/net8	vss	7.91726E-16
C2120	I0/I3922/net13	vss	7.29664E-16
C2121	I0/I3538/net13	vss	7.29758E-16
C2122	I0/I3945/net13	vss	7.20083E-16
C2123	I0/I3090/net13	vss	7.29758E-16
C2124	I0/I3561/net13	vss	7.20083E-16
C2125	I0/I3946/net13	vss	7.23918E-16
C2126	I0/I3113/net13	vss	7.20083E-16
C2127	I0/I3562/net13	vss	7.23918E-16
C2128	I0/I3935/net13	vss	7.20083E-16
C2129	I0/I3114/net13	vss	7.23918E-16
C2130	I0/I3551/net13	vss	7.20083E-16
C2131	I0/I3949/net13	vss	7.23918E-16
C2132	I0/I3103/net13	vss	7.20083E-16
C2133	I0/I3565/net13	vss	7.23918E-16
C2134	I0/I3937/net13	vss	7.20083E-16
C2135	I0/I3117/net13	vss	7.23918E-16
C2136	I0/I3553/net13	vss	7.20083E-16
C2137	I0/I3933/net13	vss	7.23918E-16
C2138	I0/I3105/net13	vss	7.20083E-16
C2139	I0/I3549/net13	vss	7.23918E-16
C2140	I0/I3939/net13	vss	7.20083E-16
C2141	I0/I3101/net13	vss	7.23918E-16
C2142	I0/I3555/net13	vss	7.20083E-16
C2143	I0/I3925/net13	vss	7.23918E-16
C2144	I0/I3107/net13	vss	7.20083E-16
C2145	I0/I3541/net13	vss	7.23918E-16
C2146	I0/I3936/net13	vss	7.20083E-16
C2147	I0/I3093/net13	vss	7.23918E-16
C2148	I0/I3552/net13	vss	7.20083E-16
C2149	I0/I3934/net13	vss	7.23918E-16
C2150	I0/I3104/net13	vss	7.20083E-16
C2151	I0/I3550/net13	vss	7.23918E-16
C2152	I0/I3928/net13	vss	7.20083E-16
C2153	I0/I3102/net13	vss	7.23918E-16
C2154	I0/I3544/net13	vss	7.20083E-16
C2155	I0/I3926/net13	vss	7.23918E-16
C2156	I0/I3096/net13	vss	7.20083E-16
C2157	I0/I3542/net13	vss	7.23918E-16
C2158	I0/I3919/net13	vss	7.20083E-16
C2159	I0/I3094/net13	vss	7.23918E-16
C2160	I0/I3535/net13	vss	7.20083E-16
C2161	I0/I3918/net13	vss	7.23918E-16
C2162	I0/I3087/net13	vss	7.20083E-16
C2163	I0/I3534/net13	vss	7.23918E-16
C2164	I0/I3940/net13	vss	7.20083E-16
C2165	I0/I3086/net13	vss	7.23918E-16
C2166	I0/I3556/net13	vss	7.20083E-16
C2167	I0/I3943/net13	vss	7.23918E-16
C2168	I0/I3108/net13	vss	7.20083E-16
C2169	I0/I3559/net13	vss	7.23918E-16
C2170	I0/I3920/net13	vss	7.20083E-16
C2171	I0/I3111/net13	vss	7.23918E-16
C2172	I0/I3536/net13	vss	7.20083E-16
C2173	I0/I3927/net13	vss	7.23918E-16
C2174	I0/I3088/net13	vss	7.20083E-16
C2175	I0/I3543/net13	vss	7.23918E-16
C2176	I0/I3941/net13	vss	7.20083E-16
C2177	I0/I3095/net13	vss	7.23918E-16
C2178	I0/I3557/net13	vss	7.20083E-16
C2179	I0/I3947/net13	vss	7.23918E-16
C2180	I0/I3109/net13	vss	7.20083E-16
C2181	I0/I3563/net13	vss	7.23918E-16
C2182	I0/I3921/net13	vss	7.20083E-16
C2183	I0/I3115/net13	vss	7.23918E-16
C2184	I0/I3537/net13	vss	7.20083E-16
C2185	I0/I3931/net13	vss	7.23918E-16
C2186	I0/I3089/net13	vss	7.20083E-16
C2187	I0/I3547/net13	vss	7.23918E-16
C2188	I0/I3930/net13	vss	7.20083E-16
C2189	I0/I3099/net13	vss	7.23918E-16
C2190	I0/I3546/net13	vss	7.20083E-16
C2191	I0/I3938/net13	vss	7.23918E-16
C2192	I0/I3098/net13	vss	7.20083E-16
C2193	I0/I3554/net13	vss	7.23918E-16
C2194	I0/I3942/net13	vss	7.20083E-16
C2195	I0/I3106/net13	vss	7.23918E-16
C2196	I0/I3558/net13	vss	7.20083E-16
C2197	I0/I3944/net13	vss	7.23918E-16
C2198	I0/I3110/net13	vss	7.20083E-16
C2199	I0/I3560/net13	vss	7.23918E-16
C2200	I0/I3929/net13	vss	7.20083E-16
C2201	I0/I3112/net13	vss	7.23918E-16
C2202	I116/net0137	vss	2.69391E-15
C2203	I0/I3545/net13	vss	7.20083E-16
C2204	I0/I3948/net13	vss	7.23918E-16
C2205	I0/I3097/net13	vss	7.20083E-16
C2206	I0/I3564/net13	vss	7.23918E-16
C2207	I0/I3923/net13	vss	7.20083E-16
C2208	I0/I3116/net13	vss	7.23918E-16
C2209	I116/net36	vss	2.5071E-15
C2210	I0/I3539/net13	vss	7.20083E-16
C2211	I0/I3924/net13	vss	7.23918E-16
C2212	I0/I3091/net13	vss	7.20083E-16
C2213	I0/I3540/net13	vss	7.23918E-16
C2214	I0/I3932/net13	vss	7.20313E-16
C2215	I0/I3092/net13	vss	7.23918E-16
C2216	I0/I3548/net13	vss	7.20313E-16
C2217	I0/I3100/net13	vss	7.20313E-16
C2218	I116/net32	vss	2.07185E-15
C2219	I1/net2224	vss	4.38252E-15
C2220	I1/net2068	vss	4.40389E-15
C2221	I1/net2212	vss	4.40979E-15
C2222	I1/net2060	vss	4.38972E-15
C2223	I1/net2152	vss	4.38594E-15
C2224	I1/net1744	vss	4.39067E-15
C2225	I1/net2140	vss	4.4022E-15
C2226	I1/net2096	vss	4.3689E-15
C2227	I0/I3922/net049	vss	9.08722E-16
C2228	I0/I3945/net049	vss	8.7222E-16
C2229	I0/I3090/net049	vss	9.09062E-16
C2230	I1/net2044	vss	4.37392E-15
C2231	I0/I3538/net049	vss	9.08793E-16
C2232	I0/I3946/net049	vss	8.95091E-16
C2233	I0/I3113/net049	vss	8.7256E-16
C2234	I0/I3561/net049	vss	8.7222E-16
C2235	I0/I3935/net049	vss	8.7222E-16
C2236	I0/I3114/net049	vss	8.95432E-16
C2237	I0/I3562/net049	vss	8.95091E-16
C2238	I0/I3949/net049	vss	8.95091E-16
C2239	I0/I3103/net049	vss	8.7256E-16
C2240	I1/net2000	vss	4.38862E-15
C2241	I0/I3551/net049	vss	8.7222E-16
C2242	I0/I3937/net049	vss	8.7222E-16
C2243	I0/I3117/net049	vss	8.95432E-16
C2244	I0/I3565/net049	vss	8.95091E-16
C2245	I0/I3933/net049	vss	8.95091E-16
C2246	I0/I3105/net049	vss	8.7256E-16
C2247	I0/I3553/net049	vss	8.7222E-16
C2248	I0/I3939/net049	vss	8.7222E-16
C2249	I0/I3101/net049	vss	8.95432E-16
C2250	I1/net1972	vss	4.38528E-15
C2251	I0/I3549/net049	vss	8.95091E-16
C2252	I0/I3925/net049	vss	8.95091E-16
C2253	I0/I3107/net049	vss	8.7256E-16
C2254	I0/I3555/net049	vss	8.7222E-16
C2255	I0/I3936/net049	vss	8.7222E-16
C2256	I0/I3093/net049	vss	8.95432E-16
C2257	I0/I3541/net049	vss	8.95091E-16
C2258	I0/I3934/net049	vss	8.95091E-16
C2259	I0/I3104/net049	vss	8.7256E-16
C2260	I1/net1944	vss	4.36783E-15
C2261	I0/I3552/net049	vss	8.7222E-16
C2262	I0/I3928/net049	vss	8.7222E-16
C2263	I0/I3102/net049	vss	8.95432E-16
C2264	I0/I3550/net049	vss	8.95091E-16
C2265	I0/I3926/net049	vss	8.95091E-16
C2266	I0/I3096/net049	vss	8.7256E-16
C2267	I0/I3544/net049	vss	8.7222E-16
C2268	I0/I3919/net049	vss	8.7222E-16
C2269	I0/I3094/net049	vss	8.95432E-16
C2270	I1/net1708	vss	4.37655E-15
C2271	I0/I3542/net049	vss	8.95091E-16
C2272	I0/I3918/net049	vss	8.95091E-16
C2273	I0/I3087/net049	vss	8.7256E-16
C2274	I0/I3535/net049	vss	8.7222E-16
C2275	I0/I3940/net049	vss	8.7222E-16
C2276	I0/I3086/net049	vss	8.95432E-16
C2277	I0/I3534/net049	vss	8.95091E-16
C2278	I0/I3943/net049	vss	8.95091E-16
C2279	I0/I3108/net049	vss	8.7256E-16
C2280	I1/net1752	vss	4.39478E-15
C2281	I0/I3556/net049	vss	8.7222E-16
C2282	I0/I3920/net049	vss	8.7222E-16
C2283	I0/I3111/net049	vss	8.95432E-16
C2284	I0/I3559/net049	vss	8.95091E-16
C2285	I0/I3927/net049	vss	8.95091E-16
C2286	I0/I3088/net049	vss	8.7256E-16
C2287	I0/I3536/net049	vss	8.7222E-16
C2288	I0/I3941/net049	vss	8.7222E-16
C2289	I0/I3095/net049	vss	8.95432E-16
C2290	I1/net1772	vss	4.3879E-15
C2291	I0/I3543/net049	vss	8.95091E-16
C2292	I0/I3947/net049	vss	8.95091E-16
C2293	I0/I3109/net049	vss	8.7256E-16
C2294	I0/I3557/net049	vss	8.7222E-16
C2295	I0/I3921/net049	vss	8.7222E-16
C2296	I0/I3115/net049	vss	8.95432E-16
C2297	I0/I3563/net049	vss	8.95091E-16
C2298	I0/I3931/net049	vss	8.95091E-16
C2299	I0/I3089/net049	vss	8.7256E-16
C2300	I1/net1904	vss	4.37359E-15
C2301	I0/I3537/net049	vss	8.7222E-16
C2302	I0/I3930/net049	vss	8.7222E-16
C2303	I0/I3099/net049	vss	8.95432E-16
C2304	I0/I3547/net049	vss	8.95091E-16
C2305	I0/I3938/net049	vss	8.95091E-16
C2306	I0/I3098/net049	vss	8.7256E-16
C2307	I0/I3546/net049	vss	8.7222E-16
C2308	I0/I3942/net049	vss	8.7222E-16
C2309	I0/I3106/net049	vss	8.95432E-16
C2310	I1/net1852	vss	4.37502E-15
C2311	I0/I3554/net049	vss	8.95091E-16
C2312	I0/I3944/net049	vss	8.95091E-16
C2313	I0/I3110/net049	vss	8.7256E-16
C2314	I0/I3558/net049	vss	8.7222E-16
C2315	I0/I3929/net049	vss	8.7222E-16
C2316	I0/I3112/net049	vss	8.95432E-16
C2317	I0/I3560/net049	vss	8.95091E-16
C2318	I0/I3948/net049	vss	8.95091E-16
C2319	I0/I3097/net049	vss	8.7256E-16
C2320	I1/net1816	vss	4.39148E-15
C2321	I0/I3545/net049	vss	8.7222E-16
C2322	I0/I3923/net049	vss	8.7222E-16
C2323	I0/I3116/net049	vss	8.95432E-16
C2324	I0/I3564/net049	vss	8.95091E-16
C2325	I0/I3924/net049	vss	8.95091E-16
C2326	I0/I3091/net049	vss	8.7256E-16
C2327	I0/I3539/net049	vss	8.7222E-16
C2328	I0/I3932/net049	vss	8.79659E-16
C2329	I0/I3092/net049	vss	8.95432E-16
C2330	I1/net1464	vss	4.4027E-15
C2331	I0/I3540/net049	vss	8.95091E-16
C2332	I0/I3100/net049	vss	8.8E-16
C2333	I0/I3548/net049	vss	8.79659E-16
C2334	I1/net1672	vss	4.3672E-15
C2335	I2/net20	vss	1.0772E-15
C2336	I5/net8	vss	7.9028E-16
C2337	I1/net1544	vss	4.37522E-15
C2338	I1/net1588	vss	4.39752E-15
C2339	I1/net1616	vss	4.40225E-15
C2340	I1/net1644	vss	4.37583E-15
C2341	I1/net1452	vss	4.37636E-15
C2342	I1/net1436	vss	4.39537E-15
C2343	I1/net1492	vss	4.40325E-15
C2344	I1/net1324	vss	4.37145E-15
C2345	I1/net1176	vss	4.37483E-15
C2346	I1/net1220	vss	4.39563E-15
C2347	I10/net8	vss	8.27156E-16
C2348	I1/net1260	vss	4.40046E-15
C2349	I2/net23	vss	5.35888E-16
C2350	I1/net1308	vss	4.4582E-15
C2351	I159/net28	vss	1.59513E-14
C2352	I116/net24	vss	3.29269E-15
C2353	I1/net1132	vss	1.56988E-15
C2354	I1/net1000	vss	1.54695E-15
C2355	I1/net1152	vss	1.54659E-15
C2356	I1/net1008	vss	1.55938E-15
C2357	I1/net560	vss	1.56293E-15
C2358	I1/net556	vss	1.54693E-15
C2359	I1/net1116	vss	1.54659E-15
C2360	I1/net1076	vss	1.5487E-15
C2361	I1/net948	vss	1.55034E-15
C2362	I1/net944	vss	1.54695E-15
C2363	I1/net908	vss	1.54659E-15
C2364	I1/net864	vss	1.54879E-15
C2365	I2/net24	vss	6.1856E-16
C2366	I1/net812	vss	1.55032E-15
C2367	I0/I3954/net13	vss	7.29927E-16
C2368	I0/I3977/net13	vss	7.19882E-16
C2369	I0/I3122/net13	vss	7.29525E-16
C2370	I1/net732	vss	1.54693E-15
C2371	I0/I3570/net13	vss	7.29664E-16
C2372	I0/I3978/net13	vss	7.23918E-16
C2373	I0/I3145/net13	vss	7.20083E-16
C2374	I0/I3593/net13	vss	7.20083E-16
C2375	I0/I3967/net13	vss	7.20083E-16
C2376	I1/net796	vss	1.54659E-15
C2377	I0/I3146/net13	vss	7.23918E-16
C2378	I0/I3594/net13	vss	7.23918E-16
C2379	I0/I3981/net13	vss	7.23918E-16
C2380	I0/I3135/net13	vss	7.20083E-16
C2381	I0/I3583/net13	vss	7.20083E-16
C2382	I0/I3969/net13	vss	7.20083E-16
C2383	I1/net788	vss	1.5487E-15
C2384	I0/I3149/net13	vss	7.23918E-16
C2385	I0/I3597/net13	vss	7.23918E-16
C2386	I0/I3965/net13	vss	7.23918E-16
C2387	I0/I3137/net13	vss	7.20083E-16
C2388	I0/I3585/net13	vss	7.20083E-16
C2389	I0/I3971/net13	vss	7.20083E-16
C2390	I1/net708	vss	1.55034E-15
C2391	I0/I3133/net13	vss	7.23918E-16
C2392	I0/I3581/net13	vss	7.23918E-16
C2393	I0/I3957/net13	vss	7.23918E-16
C2394	I0/I3139/net13	vss	7.20083E-16
C2395	I0/I3587/net13	vss	7.20083E-16
C2396	I0/I3968/net13	vss	7.20083E-16
C2397	I1/net704	vss	1.54695E-15
C2398	I0/I3125/net13	vss	7.23918E-16
C2399	I0/I3573/net13	vss	7.23918E-16
C2400	I0/I3966/net13	vss	7.23918E-16
C2401	I0/I3136/net13	vss	7.20083E-16
C2402	I0/I3584/net13	vss	7.20083E-16
C2403	I0/I3960/net13	vss	7.20083E-16
C2404	I1/net768	vss	1.54659E-15
C2405	I0/I3134/net13	vss	7.23918E-16
C2406	I0/I3582/net13	vss	7.23918E-16
C2407	I0/I3958/net13	vss	7.23918E-16
C2408	I0/I3128/net13	vss	7.20083E-16
C2409	I0/I3576/net13	vss	7.20083E-16
C2410	I0/I3951/net13	vss	7.20083E-16
C2411	I1/net600	vss	1.54879E-15
C2412	I0/I3126/net13	vss	7.23918E-16
C2413	I0/I3574/net13	vss	7.23918E-16
C2414	I0/I3950/net13	vss	7.23918E-16
C2415	I0/I3119/net13	vss	7.20083E-16
C2416	I0/I3567/net13	vss	7.20083E-16
C2417	I0/I3972/net13	vss	7.20083E-16
C2418	I0/I3118/net13	vss	7.23918E-16
C2419	I1/net452	vss	1.55032E-15
C2420	I0/I3566/net13	vss	7.23918E-16
C2421	I0/I3975/net13	vss	7.23918E-16
C2422	I0/I3140/net13	vss	7.20083E-16
C2423	I0/I3588/net13	vss	7.20083E-16
C2424	I0/I3952/net13	vss	7.20083E-16
C2425	I0/I3143/net13	vss	7.23918E-16
C2426	I1/net456	vss	1.54693E-15
C2427	I0/I3591/net13	vss	7.23918E-16
C2428	I0/I3959/net13	vss	7.23918E-16
C2429	I0/I3120/net13	vss	7.20083E-16
C2430	I0/I3568/net13	vss	7.20083E-16
C2431	I0/I3973/net13	vss	7.20083E-16
C2432	I0/I3127/net13	vss	7.23918E-16
C2433	I1/net492	vss	1.54659E-15
C2434	I0/I3575/net13	vss	7.23918E-16
C2435	I0/I3979/net13	vss	7.23918E-16
C2436	I0/I3141/net13	vss	7.20083E-16
C2437	I0/I3589/net13	vss	7.20083E-16
C2438	I0/I3953/net13	vss	7.20083E-16
C2439	I0/I3147/net13	vss	7.23918E-16
C2440	I1/net532	vss	1.54879E-15
C2441	I0/I3595/net13	vss	7.23918E-16
C2442	I0/I3963/net13	vss	7.23918E-16
C2443	I0/I3121/net13	vss	7.20083E-16
C2444	I0/I3569/net13	vss	7.20083E-16
C2445	I0/I3962/net13	vss	7.20083E-16
C2446	I0/I3131/net13	vss	7.23918E-16
C2447	I1/net352	vss	1.55034E-15
C2448	I0/I3579/net13	vss	7.23918E-16
C2449	I0/I3970/net13	vss	7.23918E-16
C2450	I0/I3130/net13	vss	7.20083E-16
C2451	I0/I3578/net13	vss	7.20083E-16
C2452	I0/I3974/net13	vss	7.20083E-16
C2453	I0/I3138/net13	vss	7.23918E-16
C2454	I1/net420	vss	1.54695E-15
C2455	I0/I3586/net13	vss	7.23918E-16
C2456	I0/I3976/net13	vss	7.23918E-16
C2457	I0/I3142/net13	vss	7.20083E-16
C2458	I0/I3590/net13	vss	7.20083E-16
C2459	I0/I3961/net13	vss	7.20083E-16
C2460	I0/I3144/net13	vss	7.23918E-16
C2461	I1/net284	vss	1.54659E-15
C2462	I0/I3592/net13	vss	7.23918E-16
C2463	I0/I3980/net13	vss	7.23918E-16
C2464	I0/I3129/net13	vss	7.20083E-16
C2465	I0/I3577/net13	vss	7.20083E-16
C2466	I0/I3955/net13	vss	7.20083E-16
C2467	I0/I3148/net13	vss	7.23918E-16
C2468	I1/net412	vss	1.54879E-15
C2469	I0/I3596/net13	vss	7.23918E-16
C2470	I0/I3956/net13	vss	7.23918E-16
C2471	I0/I3123/net13	vss	7.20083E-16
C2472	I0/I3571/net13	vss	7.20083E-16
C2473	I0/I3964/net13	vss	7.20313E-16
C2474	I0/I3124/net13	vss	7.23918E-16
C2475	I1/net72	vss	1.55032E-15
C2476	I0/I3572/net13	vss	7.23918E-16
C2477	I0/I3132/net13	vss	7.20313E-16
C2478	I0/I3580/net13	vss	7.20313E-16
C2479	I1/net76	vss	1.54693E-15
C2480	I5/net20	vss	1.07108E-15
C2481	I1/net112	vss	1.54663E-15
C2482	I1/net176	vss	1.58271E-15
C2483	I116/net0157	vss	3.2957E-15
C2484	I1/net2236	vss	1.44541E-15
C2485	I1/net2192	vss	1.50449E-15
C2486	I1/net2216	vss	1.51325E-15
C2487	I1/net2256	vss	1.55569E-15
C2488	I1/net1892	vss	1.50193E-15
C2489	I10/net20	vss	1.07168E-15
C2490	I10/net23	vss	5.28347E-16
C2491	I0/I3122/net049	vss	9.08677E-16
C2492	I5/net23	vss	5.34461E-16
C2493	I0/I3954/net049	vss	9.08677E-16
C2494	I0/I3145/net049	vss	8.7256E-16
C2495	I0/I3570/net049	vss	9.08848E-16
C2496	I0/I3977/net049	vss	8.72451E-16
C2497	I0/I3146/net049	vss	8.95432E-16
C2498	I1/net2120	vss	1.49648E-15
C2499	I0/I3593/net049	vss	8.7256E-16
C2500	I0/I3978/net049	vss	8.95432E-16
C2501	I0/I3135/net049	vss	8.7256E-16
C2502	I0/I3594/net049	vss	8.95432E-16
C2503	I0/I3967/net049	vss	8.7256E-16
C2504	I0/I3149/net049	vss	8.95432E-16
C2505	I0/I3583/net049	vss	8.7256E-16
C2506	I0/I3981/net049	vss	8.95432E-16
C2507	I0/I3137/net049	vss	8.7256E-16
C2508	I0/I3597/net049	vss	8.95432E-16
C2509	I0/I3969/net049	vss	8.7256E-16
C2510	I0/I3133/net049	vss	8.95432E-16
C2511	I1/net1396	vss	1.51325E-15
C2512	I0/I3585/net049	vss	8.7256E-16
C2513	I0/I3965/net049	vss	8.95432E-16
C2514	I0/I3139/net049	vss	8.7256E-16
C2515	I0/I3581/net049	vss	8.95432E-16
C2516	I0/I3971/net049	vss	8.7256E-16
C2517	I0/I3125/net049	vss	8.95432E-16
C2518	I0/I3587/net049	vss	8.7256E-16
C2519	I0/I3957/net049	vss	8.95432E-16
C2520	I0/I3136/net049	vss	8.7256E-16
C2521	I0/I3573/net049	vss	8.95432E-16
C2522	I0/I3968/net049	vss	8.7256E-16
C2523	I0/I3134/net049	vss	8.95432E-16
C2524	I1/net1908	vss	1.48051E-15
C2525	I0/I3584/net049	vss	8.7256E-16
C2526	I0/I3966/net049	vss	8.95432E-16
C2527	I0/I3128/net049	vss	8.7256E-16
C2528	I0/I3582/net049	vss	8.95432E-16
C2529	I0/I3960/net049	vss	8.7256E-16
C2530	I0/I3126/net049	vss	8.95432E-16
C2531	I0/I3576/net049	vss	8.7256E-16
C2532	I0/I3958/net049	vss	8.95432E-16
C2533	I0/I3119/net049	vss	8.7256E-16
C2534	I0/I3574/net049	vss	8.95432E-16
C2535	I0/I3951/net049	vss	8.7256E-16
C2536	I0/I3118/net049	vss	8.95432E-16
C2537	I1/net2032	vss	1.45167E-15
C2538	I0/I3567/net049	vss	8.7256E-16
C2539	I0/I3950/net049	vss	8.95432E-16
C2540	I0/I3140/net049	vss	8.7256E-16
C2541	I0/I3566/net049	vss	8.95432E-16
C2542	I0/I3972/net049	vss	8.7256E-16
C2543	I0/I3143/net049	vss	8.95432E-16
C2544	I0/I3588/net049	vss	8.7256E-16
C2545	I0/I3975/net049	vss	8.95432E-16
C2546	I0/I3120/net049	vss	8.7256E-16
C2547	I0/I3591/net049	vss	8.95432E-16
C2548	I0/I3952/net049	vss	8.7256E-16
C2549	I0/I3127/net049	vss	8.95432E-16
C2550	I1/net2012	vss	1.50577E-15
C2551	I0/I3568/net049	vss	8.7256E-16
C2552	I0/I3959/net049	vss	8.95432E-16
C2553	I0/I3141/net049	vss	8.7256E-16
C2554	I0/I3575/net049	vss	8.95432E-16
C2555	I0/I3973/net049	vss	8.7256E-16
C2556	I0/I3147/net049	vss	8.95432E-16
C2557	I0/I3589/net049	vss	8.7256E-16
C2558	I0/I3979/net049	vss	8.95432E-16
C2559	I0/I3121/net049	vss	8.7256E-16
C2560	I0/I3595/net049	vss	8.95432E-16
C2561	I0/I3953/net049	vss	8.7256E-16
C2562	I0/I3131/net049	vss	8.95432E-16
C2563	I1/net1984	vss	1.51325E-15
C2564	I0/I3569/net049	vss	8.7256E-16
C2565	I0/I3963/net049	vss	8.95432E-16
C2566	I0/I3130/net049	vss	8.7256E-16
C2567	I0/I3579/net049	vss	8.95432E-16
C2568	I0/I3962/net049	vss	8.7256E-16
C2569	I0/I3138/net049	vss	8.95432E-16
C2570	I0/I3578/net049	vss	8.7256E-16
C2571	I0/I3970/net049	vss	8.95432E-16
C2572	I0/I3142/net049	vss	8.7256E-16
C2573	I0/I3586/net049	vss	8.95432E-16
C2574	I0/I3974/net049	vss	8.7256E-16
C2575	I0/I3144/net049	vss	8.95432E-16
C2576	I1/net1960	vss	1.53983E-15
C2577	I0/I3590/net049	vss	8.7256E-16
C2578	I0/I3976/net049	vss	8.95432E-16
C2579	I0/I3129/net049	vss	8.7256E-16
C2580	I0/I3592/net049	vss	8.95432E-16
C2581	I0/I3961/net049	vss	8.7256E-16
C2582	I0/I3148/net049	vss	8.95432E-16
C2583	I0/I3577/net049	vss	8.7256E-16
C2584	I0/I3980/net049	vss	8.95432E-16
C2585	I0/I3123/net049	vss	8.7256E-16
C2586	I0/I3596/net049	vss	8.95432E-16
C2587	I0/I3955/net049	vss	8.7256E-16
C2588	I0/I3124/net049	vss	8.95432E-16
C2589	I1/net1484	vss	1.49274E-15
C2590	I0/I3571/net049	vss	8.7256E-16
C2591	I0/I3956/net049	vss	8.95432E-16
C2592	I0/I3132/net049	vss	8.8E-16
C2593	I0/I3572/net049	vss	8.95432E-16
C2594	I0/I3964/net049	vss	8.8E-16
C2595	I0/I3580/net049	vss	8.8E-16
C2596	I10/net24	vss	6.80049E-16
C2597	I1/net1780	vss	1.49648E-15
C2598	I5/net24	vss	6.33914E-16
C2599	I23/net7	vss	1.15941E-15
C2600	I1/net1800	vss	1.51325E-15
C2601	I1/net1716	vss	1.48051E-15
C2602	I1/net1880	vss	1.45167E-15
C2603	I1/net1352	vss	1.50577E-15
C2604	I1/net1792	vss	1.51325E-15
C2605	I1/net1840	vss	1.53983E-15
C2606	I1/net1556	vss	1.49261E-15
C2607	I1/net1576	vss	1.49648E-15
C2608	I1/net1604	vss	1.51325E-15
C2609	I1/net1628	vss	1.4806E-15
C2610	I1/net1488	vss	1.45285E-15
C2611	I1/net1496	vss	1.50577E-15
C2612	I1/net1328	vss	1.51325E-15
C2613	I1/net1420	vss	1.53983E-15
C2614	I1/net1188	vss	1.49274E-15
C2615	I1/net1208	vss	1.49648E-15
C2616	I1/net1248	vss	1.51302E-15
C2617	I0/I3602/net13	vss	7.29699E-16
C2618	I0/I3986/net13	vss	7.29837E-16
C2619	I23/net15	vss	1.17071E-15
C2620	I0/I3625/net13	vss	7.20083E-16
C2621	I0/I4009/net13	vss	7.20083E-16
C2622	I0/I3626/net13	vss	7.23918E-16
C2623	I0/I4010/net13	vss	7.23918E-16
C2624	I0/I3154/net13	vss	7.29699E-16
C2625	I0/I3615/net13	vss	7.20083E-16
C2626	I0/I3999/net13	vss	7.20083E-16
C2627	I1/net1292	vss	1.51443E-15
C2628	I0/I3177/net13	vss	7.20083E-16
C2629	I0/I3629/net13	vss	7.23918E-16
C2630	I0/I4013/net13	vss	7.23918E-16
C2631	I0/I3178/net13	vss	7.23918E-16
C2632	I0/I3617/net13	vss	7.20083E-16
C2633	I0/I4001/net13	vss	7.20083E-16
C2634	I0/I3167/net13	vss	7.20083E-16
C2635	I0/I3613/net13	vss	7.23918E-16
C2636	I0/I3997/net13	vss	7.23918E-16
C2637	I0/I3181/net13	vss	7.23918E-16
C2638	I0/I3619/net13	vss	7.20083E-16
C2639	I0/I4003/net13	vss	7.20083E-16
C2640	I0/I3169/net13	vss	7.20083E-16
C2641	I0/I3605/net13	vss	7.23918E-16
C2642	I0/I3989/net13	vss	7.23918E-16
C2643	I0/I3165/net13	vss	7.23918E-16
C2644	I116/net0149	vss	2.11431E-15
C2645	I0/I3616/net13	vss	7.20083E-16
C2646	I0/I4000/net13	vss	7.20083E-16
C2647	I0/I3171/net13	vss	7.20083E-16
C2648	I0/I3614/net13	vss	7.23918E-16
C2649	I0/I3998/net13	vss	7.23918E-16
C2650	I0/I3157/net13	vss	7.23918E-16
C2651	I1/net2184	vss	1.23989E-15
C2652	I0/I3608/net13	vss	7.20083E-16
C2653	I0/I3992/net13	vss	7.20083E-16
C2654	I0/I3168/net13	vss	7.20083E-16
C2655	I1/net2136	vss	1.23929E-15
C2656	I0/I3606/net13	vss	7.23918E-16
C2657	I0/I3990/net13	vss	7.23918E-16
C2658	I0/I3166/net13	vss	7.23918E-16
C2659	I1/net1932	vss	1.24022E-15
C2660	I0/I3599/net13	vss	7.20083E-16
C2661	I0/I3983/net13	vss	7.20083E-16
C2662	I0/I3160/net13	vss	7.20083E-16
C2663	I1/net1860	vss	1.23929E-15
C2664	I0/I3598/net13	vss	7.23918E-16
C2665	I0/I3982/net13	vss	7.23918E-16
C2666	I1/net1820	vss	1.2402E-15
C2667	I0/I3158/net13	vss	7.23918E-16
C2668	I0/I3620/net13	vss	7.20083E-16
C2669	I0/I4004/net13	vss	7.20083E-16
C2670	I1/net1656	vss	1.23931E-15
C2671	I0/I3151/net13	vss	7.20083E-16
C2672	I0/I3623/net13	vss	7.23918E-16
C2673	I0/I4007/net13	vss	7.23918E-16
C2674	I0/I3150/net13	vss	7.23918E-16
C2675	I1/net1460	vss	1.24017E-15
C2676	I0/I3600/net13	vss	7.20083E-16
C2677	I0/I3984/net13	vss	7.20083E-16
C2678	I0/I3172/net13	vss	7.20083E-16
C2679	I1/net1284	vss	1.23159E-15
C2680	I0/I3607/net13	vss	7.23918E-16
C2681	I0/I3991/net13	vss	7.23918E-16
C2682	I0/I3175/net13	vss	7.23918E-16
C2683	I0/I3621/net13	vss	7.20083E-16
C2684	I0/I4005/net13	vss	7.20083E-16
C2685	I0/I3152/net13	vss	7.20083E-16
C2686	I0/I3627/net13	vss	7.23918E-16
C2687	I0/I4011/net13	vss	7.23918E-16
C2688	I0/I3159/net13	vss	7.23918E-16
C2689	I0/I3601/net13	vss	7.20083E-16
C2690	I0/I3985/net13	vss	7.20083E-16
C2691	I0/I3173/net13	vss	7.20083E-16
C2692	I0/I3611/net13	vss	7.23918E-16
C2693	I0/I3995/net13	vss	7.23918E-16
C2694	I0/I3179/net13	vss	7.23918E-16
C2695	I0/I3610/net13	vss	7.20083E-16
C2696	I0/I3994/net13	vss	7.20083E-16
C2697	I0/I3153/net13	vss	7.20083E-16
C2698	I0/I3618/net13	vss	7.23918E-16
C2699	I0/I4002/net13	vss	7.23918E-16
C2700	I0/I3163/net13	vss	7.23918E-16
C2701	I0/I3622/net13	vss	7.20083E-16
C2702	I0/I4006/net13	vss	7.20083E-16
C2703	I0/I3162/net13	vss	7.20083E-16
C2704	I0/I3624/net13	vss	7.23918E-16
C2705	I0/I4008/net13	vss	7.23918E-16
C2706	I0/I3170/net13	vss	7.23918E-16
C2707	I0/I3609/net13	vss	7.20083E-16
C2708	I0/I3993/net13	vss	7.20083E-16
C2709	I0/I3174/net13	vss	7.20083E-16
C2710	I0/I3628/net13	vss	7.23918E-16
C2711	I0/I4012/net13	vss	7.23918E-16
C2712	I0/I3176/net13	vss	7.23918E-16
C2713	I0/I3603/net13	vss	7.20083E-16
C2714	I0/I3987/net13	vss	7.20083E-16
C2715	I0/I3161/net13	vss	7.20083E-16
C2716	I0/I3604/net13	vss	7.23918E-16
C2717	I0/I3988/net13	vss	7.23918E-16
C2718	I0/I3180/net13	vss	7.23918E-16
C2719	I0/I3612/net13	vss	7.20313E-16
C2720	I0/I3996/net13	vss	7.20313E-16
C2721	I0/I3155/net13	vss	7.20083E-16
C2722	I31/net7	vss	1.15033E-15
C2723	I0/I3156/net13	vss	7.23918E-16
C2724	I0/I3164/net13	vss	7.20313E-16
C2725	I116/net0145	vss	2.4412E-15
C2726	I1/net02030	vss	4.17428E-15
C2727	I0/I3602/net049	vss	9.09518E-16
C2728	I0/I3625/net049	vss	8.71746E-16
C2729	I0/I3986/net049	vss	9.09689E-16
C2730	I0/I3626/net049	vss	8.94618E-16
C2731	I0/I4009/net049	vss	8.71746E-16
C2732	I0/I3615/net049	vss	8.71746E-16
C2733	I0/I4010/net049	vss	8.94618E-16
C2734	I0/I3154/net049	vss	9.09518E-16
C2735	I0/I3629/net049	vss	8.94618E-16
C2736	I0/I3999/net049	vss	8.71746E-16
C2737	I0/I3177/net049	vss	8.71746E-16
C2738	I0/I3617/net049	vss	8.71746E-16
C2739	I0/I4013/net049	vss	8.94618E-16
C2740	I0/I3178/net049	vss	8.94618E-16
C2741	I0/I3613/net049	vss	8.94618E-16
C2742	I0/I4001/net049	vss	8.71746E-16
C2743	I0/I3167/net049	vss	8.71746E-16
C2744	I0/I3619/net049	vss	8.71746E-16
C2745	I0/I3997/net049	vss	8.94618E-16
C2746	I0/I3181/net049	vss	8.94618E-16
C2747	I0/I3605/net049	vss	8.94618E-16
C2748	I0/I4003/net049	vss	8.71746E-16
C2749	I0/I3169/net049	vss	8.71746E-16
C2750	I0/I3616/net049	vss	8.71746E-16
C2751	I0/I3989/net049	vss	8.94618E-16
C2752	I0/I3165/net049	vss	8.94618E-16
C2753	I0/I3614/net049	vss	8.94618E-16
C2754	I0/I4000/net049	vss	8.71746E-16
C2755	I0/I3171/net049	vss	8.71746E-16
C2756	I1/net02033	vss	9.98294E-15
C2757	I0/I3608/net049	vss	8.71746E-16
C2758	I0/I3998/net049	vss	8.94618E-16
C2759	I0/I3157/net049	vss	8.94618E-16
C2760	I1/net02041	vss	1.67737E-15
C2761	I0/I3606/net049	vss	8.94618E-16
C2762	I0/I3992/net049	vss	8.71746E-16
C2763	I0/I3168/net049	vss	8.71746E-16
C2764	I0/I3599/net049	vss	8.71746E-16
C2765	I0/I3990/net049	vss	8.94618E-16
C2766	I0/I3166/net049	vss	8.94618E-16
C2767	I0/I3598/net049	vss	8.94618E-16
C2768	I0/I3983/net049	vss	8.71746E-16
C2769	I0/I3160/net049	vss	8.71746E-16
C2770	I0/I3620/net049	vss	8.71746E-16
C2771	I0/I3982/net049	vss	8.94618E-16
C2772	I0/I3158/net049	vss	8.94618E-16
C2773	I0/I3623/net049	vss	8.94618E-16
C2774	I0/I4004/net049	vss	8.71746E-16
C2775	I0/I3151/net049	vss	8.71746E-16
C2776	I0/I3600/net049	vss	8.71746E-16
C2777	I0/I4007/net049	vss	8.94618E-16
C2778	I0/I3150/net049	vss	8.94618E-16
C2779	I0/I3607/net049	vss	8.94618E-16
C2780	I0/I3984/net049	vss	8.71746E-16
C2781	I0/I3172/net049	vss	8.71746E-16
C2782	I0/I3621/net049	vss	8.71746E-16
C2783	I0/I3991/net049	vss	8.94618E-16
C2784	I0/I3175/net049	vss	8.94618E-16
C2785	I0/I3627/net049	vss	8.94618E-16
C2786	I0/I4005/net049	vss	8.71746E-16
C2787	I0/I3152/net049	vss	8.71746E-16
C2788	I0/I3601/net049	vss	8.71746E-16
C2789	I0/I4011/net049	vss	8.94618E-16
C2790	I0/I3159/net049	vss	8.94618E-16
C2791	I1/net116	vss	7.92364E-16
C2792	I0/I3611/net049	vss	8.94618E-16
C2793	I0/I3985/net049	vss	8.71746E-16
C2794	I0/I3173/net049	vss	8.71746E-16
C2795	I1/net144	vss	7.9225E-16
C2796	I0/I3610/net049	vss	8.71746E-16
C2797	I0/I3995/net049	vss	8.94618E-16
C2798	I0/I3179/net049	vss	8.94618E-16
C2799	I1/net156	vss	7.75559E-16
C2800	I0/I3618/net049	vss	8.94618E-16
C2801	I0/I3994/net049	vss	8.71746E-16
C2802	I0/I3153/net049	vss	8.71746E-16
C2803	I0/I3622/net049	vss	8.71746E-16
C2804	I0/I4002/net049	vss	8.94618E-16
C2805	I0/I3163/net049	vss	8.94618E-16
C2806	I0/I3624/net049	vss	8.94618E-16
C2807	I0/I4006/net049	vss	8.71746E-16
C2808	I0/I3162/net049	vss	8.71746E-16
C2809	I0/I3609/net049	vss	8.71746E-16
C2810	I0/I4008/net049	vss	8.94618E-16
C2811	I0/I3170/net049	vss	8.94618E-16
C2812	I0/I3628/net049	vss	8.94618E-16
C2813	I0/I3993/net049	vss	8.71746E-16
C2814	I0/I3174/net049	vss	8.71746E-16
C2815	I0/I3603/net049	vss	8.71746E-16
C2816	I0/I4012/net049	vss	8.94618E-16
C2817	I0/I3176/net049	vss	8.94618E-16
C2818	I0/I3604/net049	vss	8.94618E-16
C2819	I0/I3987/net049	vss	8.71746E-16
C2820	I0/I3161/net049	vss	8.71746E-16
C2821	I0/I3612/net049	vss	8.79186E-16
C2822	I0/I3988/net049	vss	8.94618E-16
C2823	I0/I3180/net049	vss	8.94618E-16
C2824	I1/net336	vss	2.26389E-15
C2825	I0/I3996/net049	vss	8.79186E-16
C2826	I0/I3155/net049	vss	8.71746E-16
C2827	I26/net7	vss	1.15209E-15
C2828	I0/I3156/net049	vss	8.94618E-16
C2829	I31/net15	vss	1.18872E-15
C2830	I0/I3164/net049	vss	8.79783E-16
C2831	I1/net212	vss	1.3521E-15
C2832	I1/net320	vss	2.29834E-15
C2833	I1/net264	vss	1.37861E-15
C2834	I1/net216	vss	1.28521E-15
C2835	I1/net120	vss	1.1093E-15
C2836	I1/net328	vss	1.29667E-15
C2837	I1/net124	vss	1.11139E-15
C2838	clkout	vss	5.6779E-14
C2839	I1/net160	vss	3.63895E-15
C2840	I1/net316	vss	3.58786E-15
C2841	I1/net260	vss	2.28526E-15
C2842	I1/net516	vss	3.56571E-15
C2843	I1/net776	vss	3.58818E-15
C2844	I1/net256	vss	2.4094E-15
C2845	I1/a0bar	vss	2.12404E-14
C2846	I1/net616	vss	3.56018E-15
C2847	I1/a2bar	vss	2.06409E-14
C2848	I1/net612	vss	3.59264E-15
C2849	I1/a1	vss	2.01344E-14
C2850	I1/addr_en_b	vss	5.98287E-14
C2851	I1/net1056	vss	3.5599E-15
C2852	I1/a3	vss	3.56591E-14
C2853	I1/a3bar	vss	3.40182E-14
C2854	I1/a4	vss	3.89279E-14
C2855	I1/net880	vss	3.5881E-15
C2856	I1/a0	vss	1.68017E-14
C2857	I1/a2	vss	1.99134E-14
C2858	I1/a1bar	vss	2.03633E-14
C2859	I1/a4bar	vss	3.60534E-14
C2860	net955	vss	3.80782E-14
C2861	net954	vss	3.79851E-14
C2862	net953	vss	3.80831E-14
C2863	net951	vss	3.80302E-14
C2864	net945	vss	3.79721E-14
C2865	net943	vss	3.79252E-14
C2866	net941	vss	3.79271E-14
C2867	net939	vss	3.79053E-14
C2868	net937	vss	3.79277E-14
C2869	net935	vss	3.79382E-14
C2870	net949	vss	3.80071E-14
C2871	net947	vss	3.79642E-14
C2872	net933	vss	3.79629E-14
C2873	net929	vss	3.80146E-14
C2874	net931	vss	3.79758E-14
C2875	net927	vss	3.80452E-14
C2876	net925	vss	3.81682E-14
C2877	net924	vss	3.87171E-14
C2878	net934	vss	3.8169E-14
C2879	net926	vss	3.83128E-14
C2880	net928	vss	3.8269E-14
C2881	net930	vss	3.82465E-14
C2882	net932	vss	3.82087E-14
C2883	net936	vss	3.81562E-14
C2884	net938	vss	3.81084E-14
C2885	net940	vss	3.81227E-14
C2886	net942	vss	3.81041E-14
C2887	net944	vss	3.80713E-14
C2888	net946	vss	3.80562E-14
C2889	net948	vss	3.79985E-14
C2890	net950	vss	3.80059E-14
C2891	net952	vss	3.79866E-14
C2892	I159/net32	vss	5.73031E-15
C2893	I159/net36	vss	1.76941E-15
C2894	I33/net23	vss	1.48618E-15
C2895	BL36	vss	1.58686E-14
C2896	BL36bar	vss	2.11737E-14
C2897	p10bar	vss	6.46002E-15
C2898	BL37	vss	1.86764E-14
C2899	BL38	vss	1.89627E-14
C2900	BL39	vss	1.89799E-14
C2901	BL33	vss	1.89456E-14
C2902	BL35	vss	1.8984E-14
C2903	BL28	vss	1.89794E-14
C2904	BL29	vss	1.89728E-14
C2905	BL30	vss	1.89798E-14
C2906	BL31	vss	1.89859E-14
C2907	BL24	vss	1.89889E-14
C2908	BL25	vss	1.89685E-14
C2909	BL26	vss	1.89786E-14
C2910	BL27	vss	1.89878E-14
C2911	BL20	vss	1.89843E-14
C2912	BL21	vss	1.8969E-14
C2913	BL22	vss	1.89813E-14
C2914	BL23	vss	1.89879E-14
C2915	BL16	vss	1.89832E-14
C2916	BL17	vss	1.8947E-14
C2917	BL18	vss	1.89785E-14
C2918	BL19	vss	1.89875E-14
C2919	BL12	vss	1.89834E-14
C2920	BL13	vss	1.89671E-14
C2921	BL14	vss	1.8979E-14
C2922	BL15	vss	1.89872E-14
C2923	BL8	vss	1.89823E-14
C2924	BL9	vss	1.8973E-14
C2925	BL10	vss	1.89793E-14
C2926	BL11	vss	1.89864E-14
C2927	BL4	vss	1.89816E-14
C2928	BL5	vss	1.89683E-14
C2929	BL6	vss	1.89849E-14
C2930	BL7	vss	1.89918E-14
C2931	BL0	vss	1.89928E-14
C2932	BL1	vss	1.8978E-14
C2933	BL2	vss	1.89793E-14
C2934	BL3	vss	1.89993E-14
C2935	p10	vss	7.85874E-15
C2936	BL37bar	vss	1.89485E-14
C2937	BL38bar	vss	1.89668E-14
C2938	BL39bar	vss	1.89697E-14
C2939	BL32bar	vss	1.8972E-14
C2940	BL33bar	vss	1.89562E-14
C2941	BL34bar	vss	1.89849E-14
C2942	BL35bar	vss	1.89879E-14
C2943	BL28bar	vss	1.89713E-14
C2944	BL29bar	vss	1.89728E-14
C2945	BL30bar	vss	1.89569E-14
C2946	BL31bar	vss	1.90004E-14
C2947	BL24bar	vss	1.89806E-14
C2948	BL25bar	vss	1.89655E-14
C2949	BL26bar	vss	1.89811E-14
C2950	BL27bar	vss	1.89922E-14
C2951	BL20bar	vss	1.89728E-14
C2952	BL21bar	vss	1.89674E-14
C2953	BL22bar	vss	1.89802E-14
C2954	BL23bar	vss	1.89908E-14
C2955	BL16bar	vss	1.89714E-14
C2956	BL17bar	vss	1.89645E-14
C2957	BL18bar	vss	1.89781E-14
C2958	BL19bar	vss	1.8991E-14
C2959	BL12bar	vss	1.89718E-14
C2960	BL13bar	vss	1.89653E-14
C2961	BL14bar	vss	1.89773E-14
C2962	BL15bar	vss	1.899E-14
C2963	BL8bar	vss	1.89652E-14
C2964	BL9bar	vss	1.89654E-14
C2965	BL10bar	vss	1.89786E-14
C2966	BL11bar	vss	1.89877E-14
C2967	BL4bar	vss	1.89826E-14
C2968	BL5bar	vss	1.89693E-14
C2969	BL6bar	vss	1.89834E-14
C2970	BL7bar	vss	1.89949E-14
C2971	BL0bar	vss	1.89845E-14
C2972	BL1bar	vss	1.89426E-14
C2973	BL2bar	vss	1.89892E-14
C2974	BL3bar	vss	1.58254E-14
C2975	BL34	vss	1.89826E-14
C2976	BL32	vss	1.89804E-14
C2977	p9bar	vss	7.14698E-15
C2978	p8bar	vss	7.13043E-15
C2979	p7bar	vss	7.58044E-15
C2980	p6bar	vss	8.24237E-15
C2981	p5bar	vss	8.7195E-15
C2982	p4bar	vss	8.80901E-15
C2983	net741	vss	8.59559E-15
C2984	net256	vss	8.92836E-15
C2985	net208	vss	8.23733E-15
C2986	I32/net23	vss	1.49572E-15
C2987	I31/net23	vss	1.50576E-15
C2988	I29/net23	vss	1.50563E-15
C2989	I28/net23	vss	1.50471E-15
C2990	I27/net23	vss	1.4918E-15
C2991	I26/net23	vss	1.48343E-15
C2992	I25/net23	vss	1.48117E-15
C2993	I24/net23	vss	1.48179E-15
C2994	I23/net23	vss	1.4902E-15
C2995	p9	vss	8.35731E-15
C2996	p8	vss	8.23532E-15
C2997	p6	vss	8.8545E-15
C2998	p5	vss	9.24383E-15
C2999	p4	vss	9.53481E-15
C3000	net740	vss	9.34209E-15
C3001	net262	vss	9.65971E-15
C3002	net681	vss	2.34887E-14
C3003	net680	vss	2.0679E-14
C3004	p7	vss	8.29997E-15
C3005	I116/net0229	vss	2.5065E-15
C3006	I116/net52	vss	1.86927E-15
C3007	I116/net0309	vss	2.63176E-15
C3008	I116/net56	vss	7.0409E-15
C3009	I116/net0281	vss	2.71056E-15
C3010	I116/net60	vss	1.74406E-15
C3011	I116/net96	vss	2.75969E-15
C3012	I116/net120	vss	4.69662E-15
C3013	I116/net116	vss	2.96245E-15
C3014	I116/net0373	vss	7.47525E-15
C3015	y4bar	vss	2.72921E-14
C3016	y4	vss	2.73575E-14
C3017	y2	vss	3.13063E-14
C3018	y2bar	vss	2.90768E-14
C3019	y1bar	vss	3.07097E-14
C3020	y1	vss	2.78953E-14
C3021	y3	vss	2.49082E-14
C3022	y3bar	vss	2.26358E-14
C3023	I30/net49	vss	1.30164E-15
C3024	I30/net57	vss	3.95655E-15
C3025	I30/net61	vss	1.70299E-15
C3026	I30/net17	vss	2.40927E-15
C3027	I30/net41	vss	4.43117E-15
C3028	net220	vss	9.37625E-15
*
*
.ENDS SRAM
*
